* NGSPICE file created from heichips25_can_lehmann_fsm.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

.subckt heichips25_can_lehmann_fsm VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
X_3155_ net43 VGND VPWR net920 controller.counter2.counter_0\[2\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_3086_ net241 VGND VPWR _0109_ controller.inst_mem.mem_data\[190\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_2106_ VGND VPWR _1147_ net593 _0069_ _0328_ sg13g2_a21oi_1
X_2037_ net634 VPWR _0294_ VGND net673 net565 sg13g2_o21ai_1
XFILLER_35_461 VPWR VGND sg13g2_decap_8
X_2939_ net625 VPWR _0961_ VGND net758 net550 sg13g2_o21ai_1
Xhold351 _0187_ VPWR VGND net898 sg13g2_dlygate4sd3_1
Xhold340 _0185_ VPWR VGND net887 sg13g2_dlygate4sd3_1
Xhold362 controller.counter2.counter_1\[15\] VPWR VGND net909 sg13g2_dlygate4sd3_1
Xhold373 _0178_ VPWR VGND net920 sg13g2_dlygate4sd3_1
Xhold384 _0177_ VPWR VGND net931 sg13g2_dlygate4sd3_1
Xhold395 controller.counter2.counter_1\[12\] VPWR VGND net942 sg13g2_dlygate4sd3_1
XFILLER_41_453 VPWR VGND sg13g2_decap_8
XFILLER_36_236 VPWR VGND sg13g2_fill_1
X_2724_ net542 VPWR _0826_ VGND net893 _0773_ sg13g2_o21ai_1
X_2655_ _0771_ net448 net947 VPWR VGND sg13g2_nand2b_1
X_3207_ net79 VGND VPWR net719 controller.const_data\[22\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2586_ VGND VPWR net913 _0699_ _0706_ _1299_ sg13g2_a21oi_1
X_3138_ net105 VGND VPWR net970 controller.alu_buffer.buffer\[12\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_3069_ net275 VGND VPWR _0092_ controller.inst_mem.mem_data\[173\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
Xhold192 controller.inst_mem.mem_data\[96\] VPWR VGND net739 sg13g2_dlygate4sd3_1
Xhold170 controller.inst_mem.mem_data\[189\] VPWR VGND net717 sg13g2_dlygate4sd3_1
Xhold181 controller.extended_then_action\[1\] VPWR VGND net728 sg13g2_dlygate4sd3_1
Xfanout661 net662 net661 VPWR VGND sg13g2_buf_8
Xfanout650 net654 net650 VPWR VGND sg13g2_buf_8
X_2440_ _0583_ net485 _0582_ VPWR VGND sg13g2_nand2_1
X_2371_ VPWR VGND _0515_ _0503_ _0513_ _1069_ _0147_ _0494_ sg13g2_a221oi_1
X_2707_ net541 VPWR _0813_ VGND net924 _0773_ sg13g2_o21ai_1
X_2569_ _0692_ _0691_ net466 net455 controller.alu_buffer.buffer\[12\] VPWR VGND sg13g2_a22oi_1
X_2638_ _0753_ VPWR _0754_ VGND controller.inst_mem.mem_data\[50\] net491 sg13g2_o21ai_1
X_3120__173 VPWR VGND net173 sg13g2_tiehi
Xfanout480 _0731_ net480 VPWR VGND sg13g2_buf_8
Xfanout491 net493 net491 VPWR VGND sg13g2_buf_8
XFILLER_0_46 VPWR VGND sg13g2_fill_1
X_1940_ _1284_ _1286_ _1283_ _1287_ VPWR VGND sg13g2_nand3_1
X_1871_ _1068_ _1221_ _1222_ VPWR VGND sg13g2_nor2_1
XFILLER_6_471 VPWR VGND sg13g2_fill_2
X_2423_ _0566_ net524 controller.inst_mem.extended_word\[21\] net511 controller.inst_mem.mem_data\[173\]
+ VPWR VGND sg13g2_a22oi_1
X_2285_ VGND VPWR _0429_ _0430_ _0431_ _0428_ sg13g2_a21oi_1
X_2354_ _0499_ VPWR _0500_ VGND net777 net491 sg13g2_o21ai_1
X_3219__266 VPWR VGND net266 sg13g2_tiehi
X_3021__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_31_507 VPWR VGND sg13g2_fill_1
X_3053__307 VPWR VGND net307 sg13g2_tiehi
X_2070_ VGND VPWR _1165_ net560 _0051_ _0310_ sg13g2_a21oi_1
X_2972_ VGND VPWR _0983_ net600 _0286_ _0977_ sg13g2_a21oi_1
X_1923_ net910 net903 _1270_ _1271_ VPWR VGND sg13g2_or3_1
X_1785_ VPWR _1136_ net402 VGND sg13g2_inv_1
X_1854_ VPWR _1205_ net442 VGND sg13g2_inv_1
X_2406_ _0549_ net503 controller.inst_mem.mem_data\[199\] net507 controller.inst_mem.mem_data\[79\]
+ VPWR VGND sg13g2_a22oi_1
X_2268_ _1063_ _0410_ _1062_ _0414_ VPWR VGND _0412_ sg13g2_nand4_1
X_2337_ _0480_ _0481_ _0478_ _0483_ VPWR VGND _0482_ sg13g2_nand4_1
X_2199_ net652 VPWR _0375_ VGND net711 net599 sg13g2_o21ai_1
XFILLER_40_326 VPWR VGND sg13g2_fill_1
XFILLER_20_76 VPWR VGND sg13g2_fill_1
Xhold63 controller.const_data\[9\] VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold74 _0114_ VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold30 controller.inst_mem.mem_data\[150\] VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold52 _0103_ VPWR VGND net379 sg13g2_dlygate4sd3_1
Xhold41 controller.inst_mem.mem_data\[142\] VPWR VGND net368 sg13g2_dlygate4sd3_1
X_2985__154 VPWR VGND net154 sg13g2_tiehi
Xhold96 controller.inst_mem.mem_data\[90\] VPWR VGND net423 sg13g2_dlygate4sd3_1
Xhold85 _0059_ VPWR VGND net412 sg13g2_dlygate4sd3_1
XANTENNA_5 VPWR VGND ui_in[6] sg13g2_antennanp
X_3240_ net310 VGND VPWR net727 controller.inst_mem.mem_data\[55\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_47_492 VPWR VGND sg13g2_decap_8
X_3171_ net268 VGND VPWR net912 controller.counter2.counter_1\[2\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_1
XFILLER_39_459 VPWR VGND sg13g2_decap_8
X_2122_ VGND VPWR _1139_ net548 _0077_ _0336_ sg13g2_a21oi_1
X_2053_ net651 VPWR _0302_ VGND controller.inst_mem.mem_data\[124\] net602 sg13g2_o21ai_1
X_2955_ net655 VPWR _0969_ VGND net803 net606 sg13g2_o21ai_1
X_1768_ VPWR _1119_ net697 VGND sg13g2_inv_1
X_1837_ VPWR _1188_ net859 VGND sg13g2_inv_1
X_2886_ VGND VPWR _1026_ net582 _0243_ _0934_ sg13g2_a21oi_1
X_1906_ VGND VPWR _1257_ _1256_ _1242_ sg13g2_or2_1
X_1699_ VPWR _1050_ net713 VGND sg13g2_inv_1
XFILLER_45_407 VPWR VGND sg13g2_decap_8
XFILLER_25_153 VPWR VGND sg13g2_fill_2
Xoutput20 net20 uo_out[5] VPWR VGND sg13g2_buf_1
X_2671_ VGND VPWR _0782_ _0783_ _0178_ _0784_ sg13g2_a21oi_1
X_2740_ net911 VPWR _0838_ VGND controller.counter2.counter_1\[1\] controller.counter2.counter_1\[0\]
+ sg13g2_o21ai_1
X_3223_ net234 VGND VPWR net870 controller.inst_mem.mem_data\[38\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_3154_ net47 VGND VPWR net931 controller.counter2.counter_0\[1\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_2
X_3085_ net243 VGND VPWR net439 controller.inst_mem.mem_data\[189\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_2105_ net650 VPWR _0328_ VGND net357 net593 sg13g2_o21ai_1
X_2036_ VGND VPWR _1182_ net566 _0034_ _0293_ sg13g2_a21oi_1
X_2938_ VGND VPWR _1000_ net556 _0269_ _0960_ sg13g2_a21oi_1
Xhold363 controller.counter2.counter_1\[5\] VPWR VGND net910 sg13g2_dlygate4sd3_1
Xhold341 controller.counter2.counter_1\[6\] VPWR VGND net888 sg13g2_dlygate4sd3_1
Xhold352 controller.counter2.counter_0\[13\] VPWR VGND net899 sg13g2_dlygate4sd3_1
Xhold385 controller.counter2.counter_1\[7\] VPWR VGND net932 sg13g2_dlygate4sd3_1
Xhold374 controller.counter2.counter_1\[8\] VPWR VGND net921 sg13g2_dlygate4sd3_1
X_2869_ net658 VPWR _0926_ VGND net396 net612 sg13g2_o21ai_1
Xhold396 controller.extended_cond.opcode\[1\] VPWR VGND net943 sg13g2_dlygate4sd3_1
Xhold330 controller.inst_mem.mem_data\[38\] VPWR VGND net877 sg13g2_dlygate4sd3_1
XFILLER_45_248 VPWR VGND sg13g2_fill_2
XFILLER_41_432 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_44_281 VPWR VGND sg13g2_fill_1
X_2723_ VPWR VGND _0824_ net447 net449 net694 _0825_ net480 sg13g2_a221oi_1
X_2654_ _0767_ _0768_ _0770_ VPWR VGND sg13g2_nor2_1
X_2585_ VGND VPWR net459 _0704_ _0171_ _0705_ sg13g2_a21oi_1
X_3206_ net87 VGND VPWR _0229_ controller.const_data\[21\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3137_ net109 VGND VPWR net976 controller.alu_buffer.buffer\[11\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_2019_ net642 VPWR _1336_ VGND controller.inst_mem.mem_data\[107\] net581 sg13g2_o21ai_1
X_3068_ net277 VGND VPWR net745 controller.inst_mem.mem_data\[172\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_3107__199 VPWR VGND net199 sg13g2_tiehi
Xhold160 controller.const_data\[13\] VPWR VGND net707 sg13g2_dlygate4sd3_1
Xfanout640 net641 net640 VPWR VGND sg13g2_buf_8
Xhold171 controller.const_data\[21\] VPWR VGND net718 sg13g2_dlygate4sd3_1
Xhold182 controller.inst_mem.extended_word\[3\] VPWR VGND net729 sg13g2_dlygate4sd3_1
Xfanout651 net652 net651 VPWR VGND sg13g2_buf_8
Xhold193 controller.inst_mem.mem_data\[42\] VPWR VGND net740 sg13g2_dlygate4sd3_1
Xfanout662 net663 net662 VPWR VGND sg13g2_buf_8
XFILLER_41_251 VPWR VGND sg13g2_fill_2
XFILLER_49_340 VPWR VGND sg13g2_fill_1
X_2370_ _0494_ _0514_ _0515_ VPWR VGND sg13g2_nor2_1
X_2706_ VPWR VGND _0811_ net447 net449 net713 _0812_ net480 sg13g2_a221oi_1
XFILLER_20_479 VPWR VGND sg13g2_fill_2
X_2499_ net973 VPWR _0634_ VGND controller.alu_buffer.buffer\[6\] _1285_ sg13g2_o21ai_1
X_2568_ _1296_ net948 _0691_ VPWR VGND sg13g2_xor2_1
X_2637_ net508 controller.inst_mem.mem_data\[74\] _0752_ _0753_ VPWR VGND sg13g2_a21o_1
XFILLER_23_76 VPWR VGND sg13g2_fill_2
Xfanout470 net473 net470 VPWR VGND sg13g2_buf_8
Xfanout481 net484 net481 VPWR VGND sg13g2_buf_8
Xfanout492 net493 net492 VPWR VGND sg13g2_buf_1
X_1870_ _1221_ net533 VPWR VGND net535 sg13g2_nand2b_2
X_2995__134 VPWR VGND net134 sg13g2_tiehi
X_2422_ _0565_ controller.inst_mem.mem_data\[197\] net503 VPWR VGND sg13g2_nand2_1
X_2353_ _0496_ _0497_ _0495_ _0499_ VPWR VGND _0498_ sg13g2_nand4_1
XFILLER_37_310 VPWR VGND sg13g2_fill_2
X_2284_ _0430_ _1085_ controller.extended_cond.opcode\[1\] VPWR VGND sg13g2_nand2_1
X_3247__198 VPWR VGND net198 sg13g2_tiehi
X_1999_ net662 VPWR _1326_ VGND net421 net618 sg13g2_o21ai_1
XFILLER_19_365 VPWR VGND sg13g2_fill_1
X_1922_ controller.counter2.counter_1\[3\] controller.counter2.counter_1\[2\] controller.counter2.counter_1\[1\]
+ controller.counter2.counter_1\[0\] _1270_ VPWR VGND sg13g2_or4_1
XFILLER_34_357 VPWR VGND sg13g2_fill_1
X_2971_ net649 VPWR _0977_ VGND controller.inst_mem.mem_data\[78\] net595 sg13g2_o21ai_1
X_3236__91 VPWR VGND net91 sg13g2_tiehi
X_1853_ VPWR _1204_ net684 VGND sg13g2_inv_1
X_1784_ VPWR _1135_ net338 VGND sg13g2_inv_1
X_2336_ VGND VPWR controller.inst_mem.mem_data\[108\] net498 _0482_ net516 sg13g2_a21oi_1
X_2405_ _0548_ net495 controller.inst_mem.mem_data\[103\] net511 controller.inst_mem.mem_data\[175\]
+ VPWR VGND sg13g2_a22oi_1
X_2267_ _0410_ _0412_ _1063_ _0413_ VPWR VGND sg13g2_nand3_1
XFILLER_29_129 VPWR VGND sg13g2_fill_1
X_2198_ VGND VPWR _1101_ net603 _0115_ _0374_ sg13g2_a21oi_1
X_3189__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_48_449 VPWR VGND sg13g2_decap_8
Xhold64 _0218_ VPWR VGND net391 sg13g2_dlygate4sd3_1
Xhold86 controller.inst_mem.mem_data\[47\] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold53 controller.inst_mem.mem_data\[190\] VPWR VGND net380 sg13g2_dlygate4sd3_1
Xhold20 _0282_ VPWR VGND net347 sg13g2_dlygate4sd3_1
Xhold31 _0070_ VPWR VGND net358 sg13g2_dlygate4sd3_1
Xhold97 _0010_ VPWR VGND net424 sg13g2_dlygate4sd3_1
Xhold75 controller.inst_mem.mem_data\[160\] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold42 _0062_ VPWR VGND net369 sg13g2_dlygate4sd3_1
XANTENNA_6 VPWR VGND uio_in[0] sg13g2_antennanp
X_3196__167 VPWR VGND net167 sg13g2_tiehi
X_3170_ net272 VGND VPWR _0193_ controller.counter2.counter_1\[1\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
XFILLER_47_471 VPWR VGND sg13g2_decap_8
XFILLER_39_438 VPWR VGND sg13g2_decap_8
X_2052_ VGND VPWR _1174_ net620 _0042_ _0301_ sg13g2_a21oi_1
X_2121_ net625 VPWR _0336_ VGND net794 net548 sg13g2_o21ai_1
X_2954_ VGND VPWR _0992_ net572 _0277_ _0968_ sg13g2_a21oi_1
X_2885_ net642 VPWR _0934_ VGND net748 net582 sg13g2_o21ai_1
X_1905_ VGND VPWR _1256_ _1255_ _1249_ sg13g2_or2_1
X_1698_ VPWR _1049_ net681 VGND sg13g2_inv_1
X_1836_ VPWR _1187_ net855 VGND sg13g2_inv_1
X_1767_ VPWR _1118_ net733 VGND sg13g2_inv_1
XFILLER_1_209 VPWR VGND sg13g2_fill_2
X_2319_ _0463_ _0464_ _0465_ VPWR VGND sg13g2_and2_1
XFILLER_38_493 VPWR VGND sg13g2_decap_8
Xoutput21 net21 uo_out[6] VPWR VGND sg13g2_buf_1
X_3117__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_48_268 VPWR VGND sg13g2_fill_1
XFILLER_44_485 VPWR VGND sg13g2_decap_8
X_2670_ net540 VPWR _0784_ VGND net919 net444 sg13g2_o21ai_1
X_3153_ net51 VGND VPWR _0176_ controller.counter2.counter_0\[0\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_2
X_3222_ net242 VGND VPWR _0245_ controller.inst_mem.mem_data\[37\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2104_ VGND VPWR _1148_ net598 _0068_ _0327_ sg13g2_a21oi_1
XFILLER_35_496 VPWR VGND sg13g2_decap_8
X_2035_ net633 VPWR _0293_ VGND controller.inst_mem.mem_data\[115\] net566 sg13g2_o21ai_1
X_3084_ net245 VGND VPWR _0107_ controller.inst_mem.mem_data\[188\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_2868_ VGND VPWR _1035_ net613 _0234_ _0925_ sg13g2_a21oi_1
X_2937_ net629 VPWR _0960_ VGND controller.inst_mem.mem_data\[61\] net556 sg13g2_o21ai_1
Xhold397 controller.counter2.counter_0\[4\] VPWR VGND net944 sg13g2_dlygate4sd3_1
Xhold353 _0189_ VPWR VGND net900 sg13g2_dlygate4sd3_1
Xhold342 _0198_ VPWR VGND net889 sg13g2_dlygate4sd3_1
Xhold364 controller.counter2.counter_1\[2\] VPWR VGND net911 sg13g2_dlygate4sd3_1
X_2799_ _0884_ _0885_ _0886_ VPWR VGND sg13g2_nor2b_1
Xhold386 controller.alu_buffer.buffer\[2\] VPWR VGND net933 sg13g2_dlygate4sd3_1
Xhold375 controller.alu_buffer.buffer\[15\] VPWR VGND net922 sg13g2_dlygate4sd3_1
Xhold331 controller.extended_then_action\[5\] VPWR VGND net878 sg13g2_dlygate4sd3_1
Xhold320 controller.inst_mem.mem_data\[157\] VPWR VGND net867 sg13g2_dlygate4sd3_1
X_1819_ VPWR _1170_ net666 VGND sg13g2_inv_1
XFILLER_41_488 VPWR VGND sg13g2_decap_8
XFILLER_41_422 VPWR VGND sg13g2_fill_1
XFILLER_9_128 VPWR VGND sg13g2_fill_2
XFILLER_13_135 VPWR VGND sg13g2_fill_2
X_3234__123 VPWR VGND net123 sg13g2_tiehi
X_3245__230 VPWR VGND net230 sg13g2_tiehi
X_2722_ _0417_ net893 _0824_ VPWR VGND sg13g2_xor2_1
XFILLER_32_488 VPWR VGND sg13g2_decap_8
XFILLER_32_477 VPWR VGND sg13g2_fill_1
XFILLER_32_466 VPWR VGND sg13g2_fill_1
X_2653_ _0769_ net474 _0765_ VPWR VGND sg13g2_xnor2_1
X_2584_ net537 VPWR _0705_ VGND net956 net458 sg13g2_o21ai_1
X_3205_ net95 VGND VPWR net345 controller.const_data\[20\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3136_ net113 VGND VPWR net935 controller.alu_buffer.buffer\[10\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_3067_ net279 VGND VPWR _0090_ controller.inst_mem.mem_data\[171\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_2018_ VGND VPWR _1191_ net585 _0025_ _1335_ sg13g2_a21oi_1
XFILLER_10_105 VPWR VGND sg13g2_fill_2
Xhold172 _0230_ VPWR VGND net719 sg13g2_dlygate4sd3_1
Xfanout663 rst_n net663 VPWR VGND sg13g2_buf_8
Xfanout641 net663 net641 VPWR VGND sg13g2_buf_1
Xhold161 controller.inst_mem.mem_data\[98\] VPWR VGND net708 sg13g2_dlygate4sd3_1
Xhold150 controller.inst_mem.mem_data\[177\] VPWR VGND net697 sg13g2_dlygate4sd3_1
Xhold183 controller.inst_mem.mem_data\[111\] VPWR VGND net730 sg13g2_dlygate4sd3_1
Xfanout630 net631 net630 VPWR VGND sg13g2_buf_8
Xfanout652 net653 net652 VPWR VGND sg13g2_buf_8
Xhold194 _0251_ VPWR VGND net741 sg13g2_dlygate4sd3_1
XFILLER_37_75 VPWR VGND sg13g2_fill_1
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_37_503 VPWR VGND sg13g2_decap_4
X_2705_ _0811_ net924 _0413_ VPWR VGND sg13g2_xnor2_1
X_2636_ _0750_ _0751_ _0749_ _0752_ VPWR VGND sg13g2_nand3_1
X_2498_ VPWR VGND net967 net464 net484 net527 _0633_ net472 sg13g2_a221oi_1
X_2567_ VPWR VGND controller.alu_buffer.buffer\[21\] net461 net481 net945 _0690_ net470
+ sg13g2_a221oi_1
XFILLER_43_506 VPWR VGND sg13g2_fill_2
X_3119_ net175 VGND VPWR net354 controller.inst_mem.extended_word\[23\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
Xfanout471 net473 net471 VPWR VGND sg13g2_buf_1
Xfanout482 net484 net482 VPWR VGND sg13g2_buf_1
Xfanout460 _0596_ net460 VPWR VGND sg13g2_buf_8
Xfanout493 _1232_ net493 VPWR VGND sg13g2_buf_8
X_3199__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_34_506 VPWR VGND sg13g2_fill_2
X_2283_ _1086_ VPWR _0429_ VGND controller.extended_cond.opcode\[0\] net1 sg13g2_o21ai_1
X_2421_ _1081_ net490 _0438_ _0564_ VPWR VGND sg13g2_or3_1
X_2352_ VGND VPWR controller.inst_mem.mem_data\[176\] net503 _0498_ net517 sg13g2_a21oi_1
XFILLER_25_506 VPWR VGND sg13g2_fill_2
XFILLER_20_200 VPWR VGND sg13g2_fill_1
X_1998_ VGND VPWR _1201_ net617 _0015_ _1325_ sg13g2_a21oi_1
X_3000__124 VPWR VGND net124 sg13g2_tiehi
X_2619_ VPWR VGND controller.inst_mem.mem_data\[148\] net518 net521 controller.inst_mem.mem_data\[124\]
+ _0735_ net500 sg13g2_a221oi_1
XFILLER_28_333 VPWR VGND sg13g2_fill_2
XFILLER_1_0 VPWR VGND sg13g2_fill_2
XFILLER_19_322 VPWR VGND sg13g2_fill_2
X_1921_ net911 controller.counter2.counter_1\[1\] net892 _1269_ VPWR VGND sg13g2_nor3_1
X_1852_ VPWR _1203_ net342 VGND sg13g2_inv_1
X_2970_ VGND VPWR _0984_ net600 _0285_ _0976_ sg13g2_a21oi_1
X_1783_ VPWR _1134_ net851 VGND sg13g2_inv_1
X_2266_ controller.counter2.counter_0\[9\] controller.counter2.counter_0\[8\] _0412_
+ VPWR VGND sg13g2_nor2_1
X_2335_ _0481_ _0479_ controller.inst_mem.mem_data\[132\] net523 controller.inst_mem.extended_word\[4\]
+ VPWR VGND sg13g2_a22oi_1
X_2404_ VPWR VGND controller.inst_mem.mem_data\[151\] net518 net520 controller.inst_mem.mem_data\[127\]
+ _0547_ net499 sg13g2_a221oi_1
X_2197_ net651 VPWR _0374_ VGND controller.inst_mem.mem_data\[196\] net602 sg13g2_o21ai_1
XFILLER_48_428 VPWR VGND sg13g2_decap_8
Xhold21 controller.const_data\[15\] VPWR VGND net348 sg13g2_dlygate4sd3_1
Xhold54 _0110_ VPWR VGND net381 sg13g2_dlygate4sd3_1
Xhold10 _0088_ VPWR VGND net337 sg13g2_dlygate4sd3_1
Xhold87 controller.inst_mem.mem_data\[80\] VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold43 controller.inst_mem.mem_data\[88\] VPWR VGND net370 sg13g2_dlygate4sd3_1
Xhold76 controller.inst_mem.extended_word\[20\] VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold65 controller.inst_mem.extended_word\[19\] VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold32 controller.inst_mem.mem_data\[165\] VPWR VGND net359 sg13g2_dlygate4sd3_1
Xhold98 controller.inst_mem.mem_data\[166\] VPWR VGND net425 sg13g2_dlygate4sd3_1
XFILLER_43_188 VPWR VGND sg13g2_fill_1
XFILLER_43_177 VPWR VGND sg13g2_fill_2
XANTENNA_7 VPWR VGND uio_in[1] sg13g2_antennanp
X_2120_ VGND VPWR _1140_ net555 _0076_ _0335_ sg13g2_a21oi_1
XFILLER_47_450 VPWR VGND sg13g2_decap_8
X_2051_ net661 VPWR _0301_ VGND controller.inst_mem.mem_data\[123\] net620 sg13g2_o21ai_1
XFILLER_34_188 VPWR VGND sg13g2_fill_1
X_1835_ VPWR _1186_ net828 VGND sg13g2_inv_1
X_2884_ VGND VPWR _1027_ net583 _0242_ _0933_ sg13g2_a21oi_1
X_1904_ net514 _1022_ _1254_ _1255_ VPWR VGND sg13g2_a21o_1
X_2953_ net638 VPWR _0968_ VGND controller.inst_mem.mem_data\[69\] net572 sg13g2_o21ai_1
X_1697_ VPWR _1048_ net372 VGND sg13g2_inv_1
X_3255__254 VPWR VGND net254 sg13g2_tiehi
X_1766_ VPWR _1117_ net706 VGND sg13g2_inv_1
XFILLER_38_472 VPWR VGND sg13g2_decap_8
X_2318_ _0464_ _1019_ net515 VPWR VGND sg13g2_nand2_1
X_2249_ net653 VPWR _0400_ VGND net353 net598 sg13g2_o21ai_1
XFILLER_40_158 VPWR VGND sg13g2_fill_2
XFILLER_25_133 VPWR VGND sg13g2_fill_1
Xoutput22 net22 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_276 VPWR VGND sg13g2_fill_1
XFILLER_44_464 VPWR VGND sg13g2_decap_8
XFILLER_31_158 VPWR VGND sg13g2_fill_1
XFILLER_12_394 VPWR VGND sg13g2_fill_1
X_3221_ net250 VGND VPWR net749 controller.inst_mem.mem_data\[36\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2103_ net653 VPWR _0327_ VGND net361 net598 sg13g2_o21ai_1
X_3083_ net247 VGND VPWR net815 controller.inst_mem.mem_data\[187\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3152_ net53 VGND VPWR net918 controller.output_controller.keep\[2\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
XFILLER_35_475 VPWR VGND sg13g2_decap_8
X_3222__242 VPWR VGND net242 sg13g2_tiehi
X_2034_ VGND VPWR _1183_ net566 _0033_ _0292_ sg13g2_a21oi_1
X_2867_ net659 VPWR _0925_ VGND controller.const_data\[26\] net613 sg13g2_o21ai_1
X_2798_ net926 VPWR _0885_ VGND controller.counter2.counter_1\[12\] _1277_ sg13g2_o21ai_1
Xhold310 controller.inst_mem.mem_data\[69\] VPWR VGND net857 sg13g2_dlygate4sd3_1
X_1818_ VPWR _1169_ net798 VGND sg13g2_inv_1
X_2936_ VGND VPWR _1001_ net560 _0268_ _0959_ sg13g2_a21oi_1
Xhold365 _0194_ VPWR VGND net912 sg13g2_dlygate4sd3_1
Xhold332 controller.counter2.counter_0\[7\] VPWR VGND net879 sg13g2_dlygate4sd3_1
Xhold343 controller.counter2.counter_1\[3\] VPWR VGND net890 sg13g2_dlygate4sd3_1
Xhold354 controller.counter2.counter_1\[9\] VPWR VGND net901 sg13g2_dlygate4sd3_1
X_1749_ VPWR _1100_ net843 VGND sg13g2_inv_1
Xhold387 _0644_ VPWR VGND net934 sg13g2_dlygate4sd3_1
Xhold376 _0164_ VPWR VGND net923 sg13g2_dlygate4sd3_1
Xhold398 controller.alu_buffer.buffer\[19\] VPWR VGND net945 sg13g2_dlygate4sd3_1
Xhold321 controller.inst_mem.mem_data\[103\] VPWR VGND net868 sg13g2_dlygate4sd3_1
XFILLER_42_76 VPWR VGND sg13g2_fill_1
XFILLER_41_467 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
X_2721_ _0822_ _0823_ _0189_ VPWR VGND sg13g2_nor2_1
X_2652_ _0747_ _0765_ _0768_ VPWR VGND sg13g2_and2_1
XFILLER_8_173 VPWR VGND sg13g2_fill_1
X_3204_ net103 VGND VPWR _0227_ controller.const_data\[19\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2583_ _0702_ _0701_ _0703_ _0704_ VPWR VGND sg13g2_a21o_1
X_3135_ net117 VGND VPWR net964 controller.alu_buffer.buffer\[9\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_3066_ net281 VGND VPWR net754 controller.inst_mem.mem_data\[170\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_2017_ net643 VPWR _1335_ VGND net416 net585 sg13g2_o21ai_1
X_3028__68 VPWR VGND net68 sg13g2_tiehi
X_2919_ net646 VPWR _0951_ VGND controller.inst_mem.mem_data\[52\] net588 sg13g2_o21ai_1
Xhold140 controller.const_data\[25\] VPWR VGND net687 sg13g2_dlygate4sd3_1
Xhold162 _0018_ VPWR VGND net709 sg13g2_dlygate4sd3_1
Xhold151 _0097_ VPWR VGND net698 sg13g2_dlygate4sd3_1
XFILLER_46_504 VPWR VGND sg13g2_decap_4
Xfanout620 net621 net620 VPWR VGND sg13g2_buf_1
Xhold195 controller.inst_mem.mem_data\[123\] VPWR VGND net742 sg13g2_dlygate4sd3_1
X_3010__104 VPWR VGND net104 sg13g2_tiehi
Xhold184 _0031_ VPWR VGND net731 sg13g2_dlygate4sd3_1
Xfanout642 net645 net642 VPWR VGND sg13g2_buf_8
Xhold173 controller.inst_mem.mem_data\[33\] VPWR VGND net720 sg13g2_dlygate4sd3_1
Xfanout631 net635 net631 VPWR VGND sg13g2_buf_2
Xfanout653 net654 net653 VPWR VGND sg13g2_buf_8
X_3060__293 VPWR VGND net293 sg13g2_tiehi
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_49_320 VPWR VGND sg13g2_fill_1
X_2704_ _0809_ _0810_ _0185_ VPWR VGND sg13g2_nor2_1
X_2635_ _0751_ net525 controller.inst_mem.extended_word\[18\] net496 controller.inst_mem.mem_data\[98\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_20_459 VPWR VGND sg13g2_fill_2
X_2497_ VGND VPWR _0629_ _0631_ _0156_ _0632_ sg13g2_a21oi_1
X_2566_ VGND VPWR _0685_ _0688_ _0168_ _0689_ sg13g2_a21oi_1
X_3049_ net315 VGND VPWR net772 controller.inst_mem.mem_data\[153\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_3118_ net177 VGND VPWR _0141_ controller.inst_mem.extended_word\[22\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_23_56 VPWR VGND sg13g2_fill_2
XFILLER_46_312 VPWR VGND sg13g2_fill_2
Xfanout450 net451 net450 VPWR VGND sg13g2_buf_8
Xfanout483 net484 net483 VPWR VGND sg13g2_buf_8
Xfanout472 net473 net472 VPWR VGND sg13g2_buf_8
Xfanout461 net465 net461 VPWR VGND sg13g2_buf_8
Xfanout494 net497 net494 VPWR VGND sg13g2_buf_8
X_3242__278 VPWR VGND net278 sg13g2_tiehi
X_2420_ controller.alu_buffer.buffer\[0\] _0562_ _0563_ VPWR VGND sg13g2_nor2_1
X_2282_ net2 _0427_ _0428_ VPWR VGND sg13g2_nor2_1
X_2351_ _0497_ _0479_ controller.inst_mem.mem_data\[128\] net511 controller.inst_mem.mem_data\[152\]
+ VPWR VGND sg13g2_a22oi_1
X_1997_ net660 VPWR _1325_ VGND net739 net617 sg13g2_o21ai_1
X_2549_ VPWR VGND net952 net461 net481 controller.alu_buffer.buffer\[16\] _0675_ net470
+ sg13g2_a221oi_1
X_2618_ _0734_ net508 controller.inst_mem.mem_data\[76\] net512 controller.inst_mem.mem_data\[172\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_16_507 VPWR VGND sg13g2_fill_1
X_3127__149 VPWR VGND net149 sg13g2_tiehi
XFILLER_46_175 VPWR VGND sg13g2_fill_1
X_1851_ VPWR _1202_ net801 VGND sg13g2_inv_1
X_1920_ net17 _1267_ _1268_ VPWR VGND sg13g2_nand2_1
X_2403_ VGND VPWR _0546_ _0439_ _1079_ sg13g2_or2_1
X_1782_ VPWR _1133_ net732 VGND sg13g2_inv_1
X_2265_ _0411_ _1063_ _0410_ VPWR VGND sg13g2_nand2_1
X_2196_ VGND VPWR _1102_ net620 _0114_ _0373_ sg13g2_a21oi_1
XFILLER_27_0 VPWR VGND sg13g2_fill_1
X_2334_ _0480_ net502 controller.inst_mem.mem_data\[180\] net510 controller.inst_mem.mem_data\[156\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_48_407 VPWR VGND sg13g2_decap_8
Xhold22 _0224_ VPWR VGND net349 sg13g2_dlygate4sd3_1
Xhold11 controller.inst_mem.mem_data\[161\] VPWR VGND net338 sg13g2_dlygate4sd3_1
XFILLER_29_77 VPWR VGND sg13g2_fill_2
Xhold99 controller.inst_mem.mem_data\[57\] VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold88 _0000_ VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold44 _0008_ VPWR VGND net371 sg13g2_dlygate4sd3_1
Xhold55 controller.inst_mem.mem_data\[125\] VPWR VGND net382 sg13g2_dlygate4sd3_1
Xhold66 _0139_ VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold77 _0140_ VPWR VGND net404 sg13g2_dlygate4sd3_1
Xhold33 _0085_ VPWR VGND net360 sg13g2_dlygate4sd3_1
XANTENNA_8 VPWR VGND uio_in[2] sg13g2_antennanp
X_2050_ VGND VPWR _1175_ net621 _0041_ _0300_ sg13g2_a21oi_1
X_2952_ VGND VPWR _0993_ net572 _0276_ _0967_ sg13g2_a21oi_1
X_1834_ VPWR _1185_ net730 VGND sg13g2_inv_1
X_1765_ VPWR _1116_ net398 VGND sg13g2_inv_1
X_1903_ VGND VPWR controller.inst_mem.extended_word\[6\] net523 _1254_ _1253_ sg13g2_a21oi_1
X_2883_ net642 VPWR _0933_ VGND controller.inst_mem.mem_data\[34\] net582 sg13g2_o21ai_1
X_1696_ VPWR _1047_ net707 VGND sg13g2_inv_1
XFILLER_38_451 VPWR VGND sg13g2_decap_8
X_2179_ net634 VPWR _0365_ VGND controller.inst_mem.mem_data\[187\] net564 sg13g2_o21ai_1
X_2248_ VGND VPWR _1076_ net599 _0140_ _0399_ sg13g2_a21oi_1
X_2317_ _0460_ _0461_ _0459_ _0463_ VPWR VGND _0462_ sg13g2_nand4_1
XFILLER_31_34 VPWR VGND sg13g2_fill_1
XFILLER_48_215 VPWR VGND sg13g2_fill_1
XFILLER_44_443 VPWR VGND sg13g2_decap_8
X_3220_ net258 VGND VPWR _0243_ controller.inst_mem.mem_data\[35\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_3070__273 VPWR VGND net273 sg13g2_tiehi
X_2033_ net633 VPWR _0292_ VGND controller.inst_mem.mem_data\[114\] net566 sg13g2_o21ai_1
X_3151_ net55 VGND VPWR net941 controller.output_controller.keep\[1\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_3082_ net249 VGND VPWR net431 controller.inst_mem.mem_data\[186\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_2102_ VGND VPWR _1149_ net604 _0067_ _0326_ sg13g2_a21oi_1
XFILLER_35_454 VPWR VGND sg13g2_decap_8
X_2935_ net630 VPWR _0959_ VGND net807 net560 sg13g2_o21ai_1
Xhold344 _0195_ VPWR VGND net891 sg13g2_dlygate4sd3_1
Xhold333 _0183_ VPWR VGND net880 sg13g2_dlygate4sd3_1
X_2797_ net926 controller.counter2.counter_1\[12\] _1277_ _0884_ VPWR VGND sg13g2_nor3_1
X_2866_ VGND VPWR _1036_ net613 _0233_ _0924_ sg13g2_a21oi_1
Xhold311 controller.extended_then_action\[0\] VPWR VGND net858 sg13g2_dlygate4sd3_1
X_1748_ VPWR _1099_ net711 VGND sg13g2_inv_1
X_1817_ VPWR _1168_ net773 VGND sg13g2_inv_1
Xhold322 controller.inst_mem.mem_data\[37\] VPWR VGND net869 sg13g2_dlygate4sd3_1
Xhold300 controller.inst_mem.mem_data\[66\] VPWR VGND net847 sg13g2_dlygate4sd3_1
Xhold377 controller.counter2.counter_0\[10\] VPWR VGND net924 sg13g2_dlygate4sd3_1
Xhold355 _0201_ VPWR VGND net902 sg13g2_dlygate4sd3_1
X_1679_ VPWR _1030_ net689 VGND sg13g2_inv_1
Xhold388 _0159_ VPWR VGND net935 sg13g2_dlygate4sd3_1
X_3116__181 VPWR VGND net181 sg13g2_tiehi
Xhold366 controller.alu_buffer.buffer\[23\] VPWR VGND net913 sg13g2_dlygate4sd3_1
Xhold399 _0168_ VPWR VGND net946 sg13g2_dlygate4sd3_1
XFILLER_26_465 VPWR VGND sg13g2_fill_1
XFILLER_26_56 VPWR VGND sg13g2_fill_1
X_3240__310 VPWR VGND net310 sg13g2_tiehi
XFILLER_42_33 VPWR VGND sg13g2_fill_1
XFILLER_41_446 VPWR VGND sg13g2_decap_8
XFILLER_21_170 VPWR VGND sg13g2_fill_2
X_2720_ net542 VPWR _0823_ VGND net899 _0773_ sg13g2_o21ai_1
XFILLER_40_490 VPWR VGND sg13g2_decap_8
X_2651_ _0732_ VPWR _0767_ VGND _0747_ _0765_ sg13g2_o21ai_1
X_2582_ net950 _0562_ _0703_ VPWR VGND sg13g2_nor2_1
X_3203_ net111 VGND VPWR _0226_ controller.const_data\[18\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3134_ net121 VGND VPWR net974 controller.alu_buffer.buffer\[7\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_35_251 VPWR VGND sg13g2_fill_2
X_3065_ net283 VGND VPWR net337 controller.inst_mem.mem_data\[169\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_2016_ VGND VPWR _1192_ net592 _0024_ _1334_ sg13g2_a21oi_1
Xclkbuf_leaf_30_clk clknet_3_4__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_2918_ VGND VPWR _1010_ net588 _0259_ _0950_ sg13g2_a21oi_1
X_2849_ net640 VPWR _0916_ VGND net410 net576 sg13g2_o21ai_1
Xhold141 _0234_ VPWR VGND net688 sg13g2_dlygate4sd3_1
Xhold130 controller.inst_mem.mem_data\[82\] VPWR VGND net677 sg13g2_dlygate4sd3_1
Xhold152 controller.inst_mem.mem_data\[175\] VPWR VGND net699 sg13g2_dlygate4sd3_1
Xhold163 controller.inst_mem.extended_word\[5\] VPWR VGND net710 sg13g2_dlygate4sd3_1
Xhold174 _0242_ VPWR VGND net721 sg13g2_dlygate4sd3_1
Xhold185 controller.inst_mem.mem_data\[163\] VPWR VGND net732 sg13g2_dlygate4sd3_1
Xfanout610 net611 net610 VPWR VGND sg13g2_buf_1
Xfanout621 net622 net621 VPWR VGND sg13g2_buf_8
X_3049__315 VPWR VGND net315 sg13g2_tiehi
Xfanout643 net645 net643 VPWR VGND sg13g2_buf_8
Xfanout654 net663 net654 VPWR VGND sg13g2_buf_8
Xfanout632 net634 net632 VPWR VGND sg13g2_buf_8
Xhold196 _0043_ VPWR VGND net743 sg13g2_dlygate4sd3_1
X_3164__296 VPWR VGND net296 sg13g2_tiehi
Xclkbuf_leaf_21_clk clknet_3_6__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_12_clk clknet_3_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_2703_ net541 VPWR _0810_ VGND net886 net445 sg13g2_o21ai_1
X_2634_ _0750_ net500 controller.inst_mem.mem_data\[122\] net504 controller.inst_mem.mem_data\[194\]
+ VPWR VGND sg13g2_a22oi_1
X_2565_ net537 VPWR _0689_ VGND net945 net458 sg13g2_o21ai_1
X_2496_ net539 VPWR _0632_ VGND net527 net460 sg13g2_o21ai_1
X_3117_ net179 VGND VPWR net404 controller.inst_mem.extended_word\[21\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_3048_ net317 VGND VPWR _0071_ controller.inst_mem.mem_data\[152\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
Xfanout451 net454 net451 VPWR VGND sg13g2_buf_8
Xfanout462 net465 net462 VPWR VGND sg13g2_buf_1
Xfanout473 _0584_ net473 VPWR VGND sg13g2_buf_2
Xfanout484 _0603_ net484 VPWR VGND sg13g2_buf_8
Xfanout495 net497 net495 VPWR VGND sg13g2_buf_8
X_3015__94 VPWR VGND net94 sg13g2_tiehi
X_3030__64 VPWR VGND net64 sg13g2_tiehi
X_2281_ _0427_ controller.extended_cond.opcode\[2\] controller.extended_cond.opcode\[0\]
+ VPWR VGND sg13g2_nand2_1
X_2350_ _0496_ net495 controller.inst_mem.mem_data\[80\] net507 controller.inst_mem.mem_data\[56\]
+ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_3260__302 VPWR VGND net302 sg13g2_tiehi
X_1996_ VGND VPWR _1202_ net609 _0014_ _1324_ sg13g2_a21oi_1
X_2548_ VGND VPWR net458 _0673_ _0165_ _0674_ sg13g2_a21oi_1
X_2617_ _0733_ net525 controller.inst_mem.extended_word\[20\] net496 controller.inst_mem.mem_data\[100\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_43_316 VPWR VGND sg13g2_fill_1
X_2479_ VPWR VGND net468 net463 _0617_ net528 _0618_ net483 sg13g2_a221oi_1
Xclkload0 VPWR clkload0/Y clknet_leaf_2_clk VGND sg13g2_inv_1
XFILLER_3_445 VPWR VGND sg13g2_fill_1
XFILLER_46_198 VPWR VGND sg13g2_fill_1
XFILLER_19_346 VPWR VGND sg13g2_fill_1
XFILLER_30_500 VPWR VGND sg13g2_decap_8
X_1850_ VPWR _1201_ net821 VGND sg13g2_inv_1
X_1781_ VPWR _1132_ net714 VGND sg13g2_inv_1
X_2402_ _0537_ _0544_ _0545_ VPWR VGND sg13g2_and2_1
X_2333_ net532 net522 _0479_ VPWR VGND sg13g2_and2_1
X_2264_ net894 controller.counter2.counter_0\[5\] controller.counter2.counter_0\[4\]
+ _0410_ VGND VPWR _0407_ sg13g2_nor4_2
X_2195_ net661 VPWR _0373_ VGND controller.inst_mem.mem_data\[195\] net620 sg13g2_o21ai_1
X_3080__253 VPWR VGND net253 sg13g2_tiehi
X_1979_ net625 VPWR _1316_ VGND controller.inst_mem.mem_data\[87\] net548 sg13g2_o21ai_1
Xhold45 controller.const_data\[12\] VPWR VGND net372 sg13g2_dlygate4sd3_1
Xhold23 controller.inst_mem.mem_data\[167\] VPWR VGND net350 sg13g2_dlygate4sd3_1
Xhold56 _0045_ VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold34 controller.inst_mem.mem_data\[149\] VPWR VGND net361 sg13g2_dlygate4sd3_1
Xhold12 _0081_ VPWR VGND net339 sg13g2_dlygate4sd3_1
XFILLER_31_308 VPWR VGND sg13g2_fill_2
Xhold67 controller.inst_mem.mem_data\[191\] VPWR VGND net394 sg13g2_dlygate4sd3_1
XFILLER_28_176 VPWR VGND sg13g2_fill_2
Xhold78 controller.inst_mem.mem_data\[130\] VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold89 controller.inst_mem.mem_data\[106\] VPWR VGND net416 sg13g2_dlygate4sd3_1
XANTENNA_9 VPWR VGND uio_in[4] sg13g2_antennanp
X_3057__299 VPWR VGND net299 sg13g2_tiehi
XFILLER_47_485 VPWR VGND sg13g2_decap_8
X_1902_ _1251_ _1252_ _1250_ _1253_ VPWR VGND sg13g2_nand3_1
X_2951_ net638 VPWR _0967_ VGND net675 net572 sg13g2_o21ai_1
X_1833_ VPWR _1184_ net757 VGND sg13g2_inv_1
X_1764_ VPWR _1115_ net848 VGND sg13g2_inv_1
X_2882_ VGND VPWR _1028_ net587 _0241_ _0932_ sg13g2_a21oi_1
X_1695_ VPWR _1046_ net694 VGND sg13g2_inv_1
X_2316_ _0462_ net502 controller.inst_mem.mem_data\[185\] net510 controller.inst_mem.mem_data\[161\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_25_124 VPWR VGND sg13g2_fill_1
X_2247_ net652 VPWR _0399_ VGND controller.inst_mem.extended_word\[21\] net599 sg13g2_o21ai_1
X_2178_ VGND VPWR _1111_ net562 _0105_ _0364_ sg13g2_a21oi_1
XFILLER_5_507 VPWR VGND sg13g2_fill_1
XFILLER_44_499 VPWR VGND sg13g2_decap_8
XFILLER_44_422 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
X_3250__131 VPWR VGND net131 sg13g2_tiehi
X_3150_ net57 VGND VPWR _0173_ controller.output_controller.keep\[0\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
X_2032_ VGND VPWR _1184_ net558 _0032_ _0291_ sg13g2_a21oi_1
X_2101_ net653 VPWR _0326_ VGND controller.inst_mem.mem_data\[148\] net598 sg13g2_o21ai_1
X_3081_ net251 VGND VPWR _0104_ controller.inst_mem.mem_data\[185\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_2865_ net658 VPWR _0924_ VGND net687 net613 sg13g2_o21ai_1
X_2934_ VGND VPWR _1002_ net582 _0267_ _0958_ sg13g2_a21oi_1
Xhold356 controller.counter2.counter_1\[4\] VPWR VGND net903 sg13g2_dlygate4sd3_1
Xhold378 _0186_ VPWR VGND net925 sg13g2_dlygate4sd3_1
Xhold345 controller.counter2.counter_1\[0\] VPWR VGND net892 sg13g2_dlygate4sd3_1
X_2796_ VGND VPWR net474 _0882_ _0204_ _0883_ sg13g2_a21oi_1
X_1678_ VPWR _1029_ net873 VGND sg13g2_inv_1
Xhold367 _0172_ VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold334 controller.extended_then_action\[4\] VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold301 controller.inst_mem.mem_data\[181\] VPWR VGND net848 sg13g2_dlygate4sd3_1
X_1747_ VPWR _1098_ net755 VGND sg13g2_inv_1
X_1816_ VPWR _1167_ net340 VGND sg13g2_inv_1
Xhold312 controller.inst_mem.mem_data\[108\] VPWR VGND net859 sg13g2_dlygate4sd3_1
Xhold323 _0246_ VPWR VGND net870 sg13g2_dlygate4sd3_1
Xhold389 controller.extended_cond.opcode\[0\] VPWR VGND net936 sg13g2_dlygate4sd3_1
XFILLER_44_252 VPWR VGND sg13g2_fill_2
X_2650_ _0747_ _0765_ _0766_ VPWR VGND sg13g2_nor2_1
X_2581_ VPWR VGND net913 net456 net481 controller.alu_buffer.buffer\[21\] _0702_ net470
+ sg13g2_a221oi_1
X_3202_ net119 VGND VPWR _0225_ controller.const_data\[17\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3133_ net125 VGND VPWR _0156_ controller.alu_buffer.buffer\[6\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
X_3064_ net285 VGND VPWR _0087_ controller.inst_mem.mem_data\[168\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_2015_ net648 VPWR _1334_ VGND controller.inst_mem.mem_data\[105\] net592 sg13g2_o21ai_1
X_2848_ VGND VPWR _1045_ net578 _0224_ _0915_ sg13g2_a21oi_1
X_2917_ net646 VPWR _0950_ VGND net432 net588 sg13g2_o21ai_1
X_3192__184 VPWR VGND net184 sg13g2_tiehi
X_2779_ VGND VPWR net687 net453 _0870_ _0869_ sg13g2_a21oi_1
Xhold142 controller.const_data\[30\] VPWR VGND net689 sg13g2_dlygate4sd3_1
Xfanout622 net623 net622 VPWR VGND sg13g2_buf_2
Xfanout611 net623 net611 VPWR VGND sg13g2_buf_1
Xhold131 _0002_ VPWR VGND net678 sg13g2_dlygate4sd3_1
Xhold186 controller.inst_mem.mem_data\[178\] VPWR VGND net733 sg13g2_dlygate4sd3_1
Xfanout600 net603 net600 VPWR VGND sg13g2_buf_2
Xhold153 _0095_ VPWR VGND net700 sg13g2_dlygate4sd3_1
Xhold120 _0046_ VPWR VGND net667 sg13g2_dlygate4sd3_1
Xhold164 controller.inst_mem.mem_data\[197\] VPWR VGND net711 sg13g2_dlygate4sd3_1
Xhold175 controller.inst_mem.mem_data\[40\] VPWR VGND net722 sg13g2_dlygate4sd3_1
Xfanout633 net634 net633 VPWR VGND sg13g2_buf_8
Xhold197 controller.inst_mem.mem_data\[171\] VPWR VGND net744 sg13g2_dlygate4sd3_1
Xfanout655 net657 net655 VPWR VGND sg13g2_buf_8
Xfanout644 net645 net644 VPWR VGND sg13g2_buf_1
X_3027__70 VPWR VGND net70 sg13g2_tiehi
X_3042__40 VPWR VGND net40 sg13g2_tiehi
X_3171__268 VPWR VGND net268 sg13g2_tiehi
X_2702_ VPWR VGND _0808_ net446 net449 net390 _0809_ net480 sg13g2_a221oi_1
X_2495_ _0631_ _0630_ net469 net457 net13 VPWR VGND sg13g2_a22oi_1
X_2564_ _0688_ _0687_ net466 net455 controller.alu_buffer.buffer\[11\] VPWR VGND sg13g2_a22oi_1
X_2633_ VPWR VGND controller.inst_mem.mem_data\[146\] net518 net521 controller.inst_mem.mem_data\[170\]
+ _0749_ net512 sg13g2_a221oi_1
X_3116_ net181 VGND VPWR net393 controller.inst_mem.extended_word\[20\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_3047_ net319 VGND VPWR net358 controller.inst_mem.mem_data\[151\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
Xfanout452 net453 net452 VPWR VGND sg13g2_buf_2
Xfanout474 net475 net474 VPWR VGND sg13g2_buf_8
Xfanout463 net465 net463 VPWR VGND sg13g2_buf_8
X_3090__233 VPWR VGND net233 sg13g2_tiehi
Xfanout485 _0545_ net485 VPWR VGND sg13g2_buf_8
Xfanout496 net497 net496 VPWR VGND sg13g2_buf_2
X_2280_ net524 _0423_ _0424_ _0425_ _0426_ VPWR VGND sg13g2_nor4_1
X_3067__279 VPWR VGND net279 sg13g2_tiehi
X_2616_ _0732_ _0730_ VPWR VGND _0722_ sg13g2_nand2b_2
X_1995_ net656 VPWR _1324_ VGND controller.inst_mem.mem_data\[95\] net610 sg13g2_o21ai_1
X_2478_ _0612_ net977 _1283_ _0617_ VPWR VGND sg13g2_a21o_1
X_2547_ net537 VPWR _0674_ VGND net965 net458 sg13g2_o21ai_1
XFILLER_43_339 VPWR VGND sg13g2_fill_1
Xclkload1 clkload1/Y clknet_leaf_39_clk VPWR VGND sg13g2_inv_8
X_1780_ VPWR _1131_ net359 VGND sg13g2_inv_1
X_2401_ VGND VPWR _0475_ _0543_ _0544_ _0485_ sg13g2_a21oi_1
X_2332_ _0478_ net494 controller.inst_mem.mem_data\[84\] net506 controller.inst_mem.mem_data\[60\]
+ VPWR VGND sg13g2_a22oi_1
X_2263_ net938 controller.counter2.counter_0\[4\] _0407_ _0409_ VPWR VGND sg13g2_nor3_1
X_2194_ VGND VPWR _1103_ net619 _0113_ _0372_ sg13g2_a21oi_1
X_1978_ VGND VPWR _1211_ net557 _0005_ _1315_ sg13g2_a21oi_1
Xhold46 _0221_ VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold35 controller.inst_mem.mem_data\[122\] VPWR VGND net362 sg13g2_dlygate4sd3_1
Xhold68 _0111_ VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold79 _0050_ VPWR VGND net406 sg13g2_dlygate4sd3_1
Xhold57 controller.inst_mem.mem_data\[133\] VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold13 controller.inst_mem.mem_data\[129\] VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold24 controller.inst_mem.mem_data\[137\] VPWR VGND net351 sg13g2_dlygate4sd3_1
XFILLER_28_199 VPWR VGND sg13g2_fill_2
XFILLER_47_464 VPWR VGND sg13g2_decap_8
X_1901_ _1252_ net498 controller.inst_mem.mem_data\[110\] net506 controller.inst_mem.mem_data\[62\]
+ VPWR VGND sg13g2_a22oi_1
X_2881_ net644 VPWR _0932_ VGND net720 net587 sg13g2_o21ai_1
X_1832_ VPWR _1183_ net386 VGND sg13g2_inv_1
XFILLER_15_361 VPWR VGND sg13g2_fill_1
X_2950_ VGND VPWR _0994_ net563 _0275_ _0966_ sg13g2_a21oi_1
X_1694_ VPWR _1045_ net348 VGND sg13g2_inv_1
X_1763_ VPWR _1114_ net863 VGND sg13g2_inv_1
XFILLER_32_0 VPWR VGND sg13g2_fill_2
X_2315_ VPWR VGND controller.inst_mem.mem_data\[137\] net514 net519 controller.inst_mem.mem_data\[113\]
+ _0461_ net498 sg13g2_a221oi_1
X_2246_ VGND VPWR _1077_ net602 _0139_ _0398_ sg13g2_a21oi_1
XFILLER_38_486 VPWR VGND sg13g2_decap_8
X_2177_ net632 VPWR _0364_ VGND controller.inst_mem.mem_data\[186\] net562 sg13g2_o21ai_1
X_3167__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_44_401 VPWR VGND sg13g2_decap_8
XFILLER_44_478 VPWR VGND sg13g2_decap_8
XFILLER_16_136 VPWR VGND sg13g2_fill_1
X_3206__87 VPWR VGND net87 sg13g2_tiehi
X_3080_ net253 VGND VPWR net379 controller.inst_mem.mem_data\[184\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_2100_ VGND VPWR _1150_ net604 _0066_ _0325_ sg13g2_a21oi_1
XFILLER_35_489 VPWR VGND sg13g2_decap_8
X_2031_ net629 VPWR _0291_ VGND net386 net558 sg13g2_o21ai_1
X_2795_ net544 VPWR _0883_ VGND net942 net474 sg13g2_o21ai_1
X_2864_ VGND VPWR _1037_ net614 _0232_ _0923_ sg13g2_a21oi_1
X_1815_ VPWR _1166_ net405 VGND sg13g2_inv_1
X_2933_ net642 VPWR _0958_ VGND controller.inst_mem.mem_data\[59\] net582 sg13g2_o21ai_1
Xhold368 controller.counter2.counter_1\[1\] VPWR VGND net915 sg13g2_dlygate4sd3_1
Xhold346 controller.counter2.counter_0\[14\] VPWR VGND net893 sg13g2_dlygate4sd3_1
Xhold379 controller.counter2.counter_1\[13\] VPWR VGND net926 sg13g2_dlygate4sd3_1
Xhold357 controller.counter2.counter_1\[14\] VPWR VGND net904 sg13g2_dlygate4sd3_1
Xhold335 controller.extended_then_action\[3\] VPWR VGND net882 sg13g2_dlygate4sd3_1
Xhold302 _0101_ VPWR VGND net849 sg13g2_dlygate4sd3_1
X_1746_ VPWR _1097_ net829 VGND sg13g2_inv_1
Xhold324 controller.inst_mem.mem_data\[159\] VPWR VGND net871 sg13g2_dlygate4sd3_1
X_1677_ VPWR _1028_ net777 VGND sg13g2_inv_1
Xhold313 controller.inst_mem.mem_data\[101\] VPWR VGND net860 sg13g2_dlygate4sd3_1
X_2229_ net638 VPWR _0390_ VGND net858 net575 sg13g2_o21ai_1
X_3123__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_12_183 VPWR VGND sg13g2_fill_2
XFILLER_16_91 VPWR VGND sg13g2_fill_1
X_2580_ _0701_ net467 _0700_ VPWR VGND sg13g2_nand2_1
X_3201_ net127 VGND VPWR net349 controller.const_data\[16\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3132_ net129 VGND VPWR net962 controller.alu_buffer.buffer\[5\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_3063_ net287 VGND VPWR _0086_ controller.inst_mem.mem_data\[167\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_2981__162 VPWR VGND net162 sg13g2_tiehi
X_2014_ VGND VPWR _1193_ net597 _0023_ _1333_ sg13g2_a21oi_1
X_2847_ net640 VPWR _0915_ VGND controller.const_data\[16\] net578 sg13g2_o21ai_1
X_2778_ net453 _0868_ _0869_ VPWR VGND sg13g2_nor2_1
X_2916_ VGND VPWR _1011_ net608 _0258_ _0949_ sg13g2_a21oi_1
X_3077__259 VPWR VGND net259 sg13g2_tiehi
Xhold110 _0067_ VPWR VGND net437 sg13g2_dlygate4sd3_1
Xfanout612 net614 net612 VPWR VGND sg13g2_buf_8
Xfanout623 net624 net623 VPWR VGND sg13g2_buf_2
Xhold143 _0239_ VPWR VGND net690 sg13g2_dlygate4sd3_1
Xhold187 controller.inst_mem.mem_data\[72\] VPWR VGND net734 sg13g2_dlygate4sd3_1
Xfanout656 net657 net656 VPWR VGND sg13g2_buf_8
X_1729_ VPWR _1080_ net881 VGND sg13g2_inv_1
Xhold154 controller.inst_mem.extended_word\[6\] VPWR VGND net701 sg13g2_dlygate4sd3_1
Xhold121 controller.inst_mem.mem_data\[135\] VPWR VGND net668 sg13g2_dlygate4sd3_1
Xfanout645 net654 net645 VPWR VGND sg13g2_buf_8
Xhold165 _0117_ VPWR VGND net712 sg13g2_dlygate4sd3_1
Xhold176 _0249_ VPWR VGND net723 sg13g2_dlygate4sd3_1
Xfanout634 net635 net634 VPWR VGND sg13g2_buf_8
Xhold198 _0091_ VPWR VGND net745 sg13g2_dlygate4sd3_1
Xfanout601 net602 net601 VPWR VGND sg13g2_buf_8
Xhold132 controller.inst_mem.mem_data\[145\] VPWR VGND net679 sg13g2_dlygate4sd3_1
XFILLER_41_245 VPWR VGND sg13g2_fill_1
XFILLER_41_223 VPWR VGND sg13g2_fill_2
XFILLER_14_415 VPWR VGND sg13g2_fill_1
XFILLER_14_426 VPWR VGND sg13g2_fill_1
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_37_507 VPWR VGND sg13g2_fill_1
XFILLER_1_374 VPWR VGND sg13g2_fill_2
X_3137__109 VPWR VGND net109 sg13g2_tiehi
X_2701_ _0808_ _0413_ _0807_ VPWR VGND sg13g2_nand2_1
X_2632_ _0739_ net487 _0746_ _0748_ VPWR VGND sg13g2_a21o_2
X_2494_ _0630_ net527 _1285_ VPWR VGND sg13g2_xnor2_1
X_2563_ _0687_ _0686_ _1296_ VPWR VGND sg13g2_nand2b_1
X_3046_ net321 VGND VPWR _0069_ controller.inst_mem.mem_data\[150\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_3115_ net183 VGND VPWR net365 controller.inst_mem.extended_word\[19\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
Xfanout464 net465 net464 VPWR VGND sg13g2_buf_1
Xfanout453 net454 net453 VPWR VGND sg13g2_buf_8
Xfanout475 _0748_ net475 VPWR VGND sg13g2_buf_8
Xfanout486 _0474_ net486 VPWR VGND sg13g2_buf_8
Xfanout497 _1227_ net497 VPWR VGND sg13g2_buf_8
XFILLER_19_507 VPWR VGND sg13g2_fill_1
X_3214__306 VPWR VGND net306 sg13g2_tiehi
XFILLER_6_488 VPWR VGND sg13g2_fill_2
X_1994_ VGND VPWR _1203_ net607 _0013_ _1323_ sg13g2_a21oi_1
X_2615_ _0722_ _0730_ _0731_ VPWR VGND sg13g2_nor2b_1
X_2477_ VGND VPWR _0611_ _0615_ _0152_ _0616_ sg13g2_a21oi_1
X_2546_ _0672_ _0671_ _0668_ _0673_ VPWR VGND sg13g2_a21o_1
X_3029_ net66 VGND VPWR _0052_ controller.inst_mem.mem_data\[133\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
Xclkload2 clknet_leaf_34_clk clkload2/Y VPWR VGND sg13g2_inv_4
X_2400_ _0542_ VPWR _0543_ VGND controller.inst_mem.mem_data\[48\] net492 sg13g2_o21ai_1
X_3251__99 VPWR VGND net99 sg13g2_tiehi
X_2262_ net944 _0407_ _0408_ VPWR VGND sg13g2_nor2_1
X_2331_ _0477_ net486 _0476_ VPWR VGND sg13g2_nand2_1
XFILLER_37_156 VPWR VGND sg13g2_fill_2
X_2193_ net661 VPWR _0372_ VGND net400 net619 sg13g2_o21ai_1
X_1977_ net628 VPWR _1315_ VGND net784 net550 sg13g2_o21ai_1
X_2529_ net538 VPWR _0659_ VGND net954 net459 sg13g2_o21ai_1
XFILLER_20_38 VPWR VGND sg13g2_fill_2
Xhold69 controller.const_data\[27\] VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold36 _0042_ VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold14 _0049_ VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold58 _0053_ VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold47 controller.inst_mem.mem_data\[65\] VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold25 _0057_ VPWR VGND net352 sg13g2_dlygate4sd3_1
XFILLER_47_443 VPWR VGND sg13g2_decap_8
X_3209__63 VPWR VGND net63 sg13g2_tiehi
X_1900_ _1251_ net502 controller.inst_mem.mem_data\[182\] net510 controller.inst_mem.mem_data\[158\]
+ VPWR VGND sg13g2_a22oi_1
X_1831_ VPWR _1182_ net763 VGND sg13g2_inv_1
X_3105__203 VPWR VGND net203 sg13g2_tiehi
X_2880_ VGND VPWR _1029_ net590 _0240_ _0931_ sg13g2_a21oi_1
X_1693_ VPWR _1044_ net418 VGND sg13g2_inv_1
X_1762_ VPWR _1113_ net378 VGND sg13g2_inv_1
XFILLER_38_465 VPWR VGND sg13g2_decap_8
X_2176_ VGND VPWR _1112_ net551 _0104_ _0363_ sg13g2_a21oi_1
X_2314_ _0460_ net523 controller.extended_cond.opcode\[0\] net506 controller.inst_mem.mem_data\[65\]
+ VPWR VGND sg13g2_a22oi_1
X_2245_ net651 VPWR _0398_ VGND controller.inst_mem.extended_word\[20\] net602 sg13g2_o21ai_1
X_3006__112 VPWR VGND net112 sg13g2_tiehi
X_3195__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_33_192 VPWR VGND sg13g2_fill_2
X_2991__142 VPWR VGND net142 sg13g2_tiehi
Xoutput15 net15 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_44_457 VPWR VGND sg13g2_decap_8
X_3087__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_12_354 VPWR VGND sg13g2_fill_1
X_3174__256 VPWR VGND net256 sg13g2_tiehi
X_2030_ VGND VPWR _1185_ net550 _0031_ _0290_ sg13g2_a21oi_1
XFILLER_35_468 VPWR VGND sg13g2_decap_8
X_2932_ VGND VPWR _1003_ net591 _0266_ _0957_ sg13g2_a21oi_1
X_2863_ net659 VPWR _0923_ VGND net811 net613 sg13g2_o21ai_1
X_2794_ VGND VPWR net822 net450 _0882_ _0881_ sg13g2_a21oi_1
X_1814_ VPWR _1165_ net831 VGND sg13g2_inv_1
XFILLER_7_61 VPWR VGND sg13g2_fill_2
X_1745_ VPWR _1096_ net844 VGND sg13g2_inv_1
Xhold369 controller.counter2.counter_0\[12\] VPWR VGND net916 sg13g2_dlygate4sd3_1
Xhold347 controller.counter2.counter_0\[6\] VPWR VGND net894 sg13g2_dlygate4sd3_1
Xhold358 _0206_ VPWR VGND net905 sg13g2_dlygate4sd3_1
Xhold336 controller.counter2.counter_1\[11\] VPWR VGND net883 sg13g2_dlygate4sd3_1
X_1676_ VPWR _1027_ net720 VGND sg13g2_inv_1
Xhold303 controller.inst_mem.mem_data\[176\] VPWR VGND net850 sg13g2_dlygate4sd3_1
Xhold314 _0021_ VPWR VGND net861 sg13g2_dlygate4sd3_1
Xhold325 controller.inst_mem.mem_data\[55\] VPWR VGND net872 sg13g2_dlygate4sd3_1
X_2228_ VGND VPWR _1086_ net575 _0130_ _0389_ sg13g2_a21oi_1
X_2159_ net648 VPWR _0355_ VGND net697 net592 sg13g2_o21ai_1
Xclkbuf_leaf_33_clk clknet_3_1__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_3130__137 VPWR VGND net137 sg13g2_tiehi
Xclkbuf_leaf_24_clk clknet_3_5__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
X_3200_ net135 VGND VPWR _0223_ controller.const_data\[15\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_4_361 VPWR VGND sg13g2_fill_1
X_3131_ net133 VGND VPWR net981 controller.alu_buffer.buffer\[4\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_2013_ net649 VPWR _1333_ VGND net388 net597 sg13g2_o21ai_1
X_3062_ net289 VGND VPWR net360 controller.inst_mem.mem_data\[166\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_15_clk clknet_3_6__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_2915_ net656 VPWR _0949_ VGND net434 net608 sg13g2_o21ai_1
X_2846_ VGND VPWR _1046_ net577 _0223_ _0914_ sg13g2_a21oi_1
X_2777_ _1274_ _0867_ _0868_ VPWR VGND sg13g2_nor2b_1
Xhold122 controller.inst_mem.mem_data\[71\] VPWR VGND net669 sg13g2_dlygate4sd3_1
XFILLER_31_493 VPWR VGND sg13g2_decap_8
X_1728_ _1079_ net878 VPWR VGND sg13g2_inv_2
Xhold100 _0266_ VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold144 controller.inst_mem.mem_data\[79\] VPWR VGND net691 sg13g2_dlygate4sd3_1
Xhold133 _0065_ VPWR VGND net680 sg13g2_dlygate4sd3_1
Xhold111 controller.inst_mem.mem_data\[188\] VPWR VGND net438 sg13g2_dlygate4sd3_1
Xhold166 controller.const_data\[10\] VPWR VGND net713 sg13g2_dlygate4sd3_1
Xfanout624 _1309_ net624 VPWR VGND sg13g2_buf_8
Xfanout613 net614 net613 VPWR VGND sg13g2_buf_8
Xfanout657 net659 net657 VPWR VGND sg13g2_buf_8
X_1659_ VPWR _1010_ net434 VGND sg13g2_inv_1
Xhold177 controller.inst_mem.mem_data\[84\] VPWR VGND net724 sg13g2_dlygate4sd3_1
Xhold155 _0126_ VPWR VGND net702 sg13g2_dlygate4sd3_1
Xhold188 controller.inst_mem.mem_data\[148\] VPWR VGND net735 sg13g2_dlygate4sd3_1
Xfanout635 net663 net635 VPWR VGND sg13g2_buf_8
Xfanout646 net654 net646 VPWR VGND sg13g2_buf_8
Xhold199 controller.inst_mem.mem_data\[124\] VPWR VGND net746 sg13g2_dlygate4sd3_1
Xfanout602 net603 net602 VPWR VGND sg13g2_buf_8
X_3201__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_49_368 VPWR VGND sg13g2_decap_8
X_2700_ net886 VPWR _0807_ VGND controller.counter2.counter_0\[8\] _0411_ sg13g2_o21ai_1
X_2631_ VGND VPWR _0746_ _0747_ _0739_ net487 sg13g2_a21oi_2
X_2562_ _0686_ net945 _0680_ VPWR VGND sg13g2_nand2b_1
X_2493_ VPWR VGND net973 net464 net483 net980 _0629_ net472 sg13g2_a221oi_1
X_3113__187 VPWR VGND net187 sg13g2_tiehi
Xclkbuf_leaf_4_clk clknet_3_6__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_3114_ net185 VGND VPWR _0137_ controller.inst_mem.extended_word\[18\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_3045_ net323 VGND VPWR _0068_ controller.inst_mem.mem_data\[149\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_2829_ net636 VPWR _0906_ VGND controller.const_data\[7\] net569 sg13g2_o21ai_1
Xfanout454 _0830_ net454 VPWR VGND sg13g2_buf_8
Xfanout476 net477 net476 VPWR VGND sg13g2_buf_8
Xfanout465 _0595_ net465 VPWR VGND sg13g2_buf_2
Xfanout487 _0474_ net487 VPWR VGND sg13g2_buf_1
Xfanout498 net501 net498 VPWR VGND sg13g2_buf_8
XFILLER_33_500 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_45_393 VPWR VGND sg13g2_decap_8
X_1993_ net655 VPWR _1323_ VGND controller.inst_mem.mem_data\[94\] net607 sg13g2_o21ai_1
X_2614_ VGND VPWR _0475_ _0729_ _0730_ _0485_ sg13g2_a21oi_1
X_2545_ VPWR VGND net958 net455 net481 net922 _0672_ net470 sg13g2_a221oi_1
X_2476_ net539 VPWR _0616_ VGND net529 net460 sg13g2_o21ai_1
X_3028_ net68 VGND VPWR _0051_ controller.inst_mem.mem_data\[132\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
Xclkload3 clkload3/Y clknet_leaf_6_clk VPWR VGND sg13g2_inv_8
XFILLER_3_404 VPWR VGND sg13g2_fill_1
XFILLER_42_352 VPWR VGND sg13g2_fill_2
X_3066__281 VPWR VGND net281 sg13g2_tiehi
X_3097__219 VPWR VGND net219 sg13g2_tiehi
X_2261_ controller.counter2.counter_0\[3\] controller.counter2.counter_0\[2\] controller.counter2.counter_0\[1\]
+ controller.counter2.counter_0\[0\] _0407_ VPWR VGND sg13g2_or4_1
X_2192_ VGND VPWR _1104_ net618 _0112_ _0371_ sg13g2_a21oi_1
X_2330_ VGND VPWR net535 net488 _0476_ _0440_ sg13g2_a21oi_1
X_1976_ VGND VPWR _1212_ net555 _0004_ _1314_ sg13g2_a21oi_1
X_2528_ _0658_ _0657_ net467 net456 controller.alu_buffer.buffer\[5\] VPWR VGND sg13g2_a22oi_1
X_2978__168 VPWR VGND net168 sg13g2_tiehi
X_2459_ net538 VPWR _0602_ VGND net967 _0601_ sg13g2_o21ai_1
Xhold37 controller.inst_mem.extended_word\[18\] VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold15 controller.inst_mem.mem_data\[93\] VPWR VGND net342 sg13g2_dlygate4sd3_1
Xhold59 controller.inst_mem.mem_data\[113\] VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold26 controller.inst_mem.extended_word\[22\] VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold48 _0274_ VPWR VGND net375 sg13g2_dlygate4sd3_1
X_3126__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_47_422 VPWR VGND sg13g2_decap_8
XFILLER_3_267 VPWR VGND sg13g2_fill_2
XFILLER_47_499 VPWR VGND sg13g2_decap_8
XFILLER_19_70 VPWR VGND sg13g2_fill_2
XFILLER_19_81 VPWR VGND sg13g2_fill_2
X_1761_ VPWR _1112_ net846 VGND sg13g2_inv_1
X_1830_ VPWR _1181_ net819 VGND sg13g2_inv_1
X_1692_ VPWR _1043_ net410 VGND sg13g2_inv_1
X_2313_ _0459_ controller.inst_mem.mem_data\[89\] net494 VPWR VGND sg13g2_nand2_1
XFILLER_38_444 VPWR VGND sg13g2_decap_8
X_2175_ net626 VPWR _0363_ VGND net430 net551 sg13g2_o21ai_1
XFILLER_18_0 VPWR VGND sg13g2_fill_1
X_2244_ VGND VPWR _1078_ net602 _0138_ _0397_ sg13g2_a21oi_1
X_1959_ net20 _1303_ _1304_ VPWR VGND sg13g2_nand2_2
Xoutput16 net16 uo_out[1] VPWR VGND sg13g2_buf_1
X_3151__55 VPWR VGND net55 sg13g2_tiehi
XFILLER_44_436 VPWR VGND sg13g2_decap_8
X_3204__103 VPWR VGND net103 sg13g2_tiehi
X_3215__298 VPWR VGND net298 sg13g2_tiehi
X_3181__228 VPWR VGND net228 sg13g2_tiehi
XFILLER_35_447 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_2931_ net644 VPWR _0957_ VGND controller.inst_mem.mem_data\[58\] net583 sg13g2_o21ai_1
X_2862_ VGND VPWR _1038_ net613 _0231_ _0922_ sg13g2_a21oi_1
X_2793_ net450 _0880_ _0881_ VPWR VGND sg13g2_nor2_1
Xhold326 controller.const_data\[31\] VPWR VGND net873 sg13g2_dlygate4sd3_1
X_1813_ VPWR _1164_ net692 VGND sg13g2_inv_1
X_1744_ VPWR _1095_ net854 VGND sg13g2_inv_1
Xhold315 controller.inst_mem.mem_data\[63\] VPWR VGND net862 sg13g2_dlygate4sd3_1
Xhold304 controller.inst_mem.mem_data\[162\] VPWR VGND net851 sg13g2_dlygate4sd3_1
Xhold359 controller.counter2.counter_0\[15\] VPWR VGND net906 sg13g2_dlygate4sd3_1
Xhold348 _0182_ VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold337 _0203_ VPWR VGND net884 sg13g2_dlygate4sd3_1
X_1675_ VPWR _1026_ net800 VGND sg13g2_inv_1
XFILLER_41_406 VPWR VGND sg13g2_fill_2
X_2227_ net639 VPWR _0389_ VGND net885 net575 sg13g2_o21ai_1
X_2158_ VGND VPWR _1121_ net597 _0095_ _0354_ sg13g2_a21oi_1
X_2089_ net646 VPWR _0320_ VGND controller.inst_mem.mem_data\[142\] net590 sg13g2_o21ai_1
XFILLER_41_439 VPWR VGND sg13g2_decap_8
XFILLER_13_119 VPWR VGND sg13g2_fill_2
XFILLER_32_417 VPWR VGND sg13g2_fill_1
XFILLER_40_483 VPWR VGND sg13g2_decap_8
X_3130_ net137 VGND VPWR _0153_ controller.alu_buffer.buffer\[3\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_2
X_2012_ VGND VPWR _1194_ net595 _0022_ _1332_ sg13g2_a21oi_1
X_3061_ net291 VGND VPWR _0084_ controller.inst_mem.mem_data\[165\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_2845_ net640 VPWR _0914_ VGND net348 net577 sg13g2_o21ai_1
X_2914_ VGND VPWR _1012_ net609 _0257_ _0948_ sg13g2_a21oi_1
Xhold134 controller.const_data\[11\] VPWR VGND net681 sg13g2_dlygate4sd3_1
X_2776_ net901 VPWR _0867_ VGND controller.counter2.counter_1\[8\] _1273_ sg13g2_o21ai_1
Xhold123 _0280_ VPWR VGND net670 sg13g2_dlygate4sd3_1
X_1727_ VPWR _1078_ net364 VGND sg13g2_inv_1
Xhold112 _0108_ VPWR VGND net439 sg13g2_dlygate4sd3_1
Xhold156 controller.inst_mem.mem_data\[155\] VPWR VGND net703 sg13g2_dlygate4sd3_1
Xhold101 controller.inst_mem.mem_data\[134\] VPWR VGND net428 sg13g2_dlygate4sd3_1
Xhold145 controller.inst_mem.mem_data\[132\] VPWR VGND net692 sg13g2_dlygate4sd3_1
X_1658_ VPWR _1009_ net432 VGND sg13g2_inv_1
Xhold167 controller.inst_mem.mem_data\[164\] VPWR VGND net714 sg13g2_dlygate4sd3_1
Xfanout636 net637 net636 VPWR VGND sg13g2_buf_8
Xhold189 controller.const_data\[20\] VPWR VGND net736 sg13g2_dlygate4sd3_1
Xfanout658 net659 net658 VPWR VGND sg13g2_buf_8
Xfanout614 net623 net614 VPWR VGND sg13g2_buf_8
X_3259_ net83 VGND VPWR net347 controller.inst_mem.mem_data\[74\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
Xfanout647 net654 net647 VPWR VGND sg13g2_buf_1
Xhold178 _0004_ VPWR VGND net725 sg13g2_dlygate4sd3_1
Xfanout625 net626 net625 VPWR VGND sg13g2_buf_8
Xfanout603 net604 net603 VPWR VGND sg13g2_buf_8
XFILLER_41_225 VPWR VGND sg13g2_fill_1
XFILLER_17_200 VPWR VGND sg13g2_fill_2
XFILLER_13_450 VPWR VGND sg13g2_fill_2
X_2492_ VPWR VGND _0628_ _0503_ _0627_ _1066_ _0155_ net464 sg13g2_a221oi_1
X_2630_ _0486_ VPWR _0746_ VGND net487 _0745_ sg13g2_o21ai_1
X_2561_ VPWR VGND controller.alu_buffer.buffer\[20\] net461 net481 controller.alu_buffer.buffer\[18\]
+ _0685_ net470 sg13g2_a221oi_1
X_3076__261 VPWR VGND net261 sg13g2_tiehi
X_3113_ net187 VGND VPWR _0136_ controller.extended_then_action\[5\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_3044_ net325 VGND VPWR net437 controller.inst_mem.mem_data\[148\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_2828_ VGND VPWR _1055_ net569 _0214_ _0905_ sg13g2_a21oi_1
X_3024__76 VPWR VGND net76 sg13g2_tiehi
X_2759_ net544 VPWR _0854_ VGND net910 net476 sg13g2_o21ai_1
Xfanout444 net445 net444 VPWR VGND sg13g2_buf_8
Xfanout477 net478 net477 VPWR VGND sg13g2_buf_2
Xfanout455 net456 net455 VPWR VGND sg13g2_buf_8
Xfanout488 _0439_ net488 VPWR VGND sg13g2_buf_8
Xfanout466 net467 net466 VPWR VGND sg13g2_buf_8
X_2988__148 VPWR VGND net148 sg13g2_tiehi
Xfanout499 net501 net499 VPWR VGND sg13g2_buf_8
Xclkload10 clknet_leaf_18_clk clkload10/X VPWR VGND sg13g2_buf_8
X_1992_ VGND VPWR _1204_ net572 _0012_ _1322_ sg13g2_a21oi_1
X_2475_ _0615_ _0614_ net468 net457 net9 VPWR VGND sg13g2_a22oi_1
X_2613_ VPWR _0729_ _0728_ VGND sg13g2_inv_1
X_2544_ net466 VPWR _0671_ VGND _0669_ _0670_ sg13g2_o21ai_1
XFILLER_36_361 VPWR VGND sg13g2_fill_2
X_3027_ net70 VGND VPWR net406 controller.inst_mem.mem_data\[131\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_3241__294 VPWR VGND net294 sg13g2_tiehi
XFILLER_11_239 VPWR VGND sg13g2_fill_1
Xclkload4 VPWR clkload4/Y clknet_leaf_7_clk VGND sg13g2_inv_1
X_3177__244 VPWR VGND net244 sg13g2_tiehi
X_3218__274 VPWR VGND net274 sg13g2_tiehi
X_2191_ net662 VPWR _0371_ VGND net682 net621 sg13g2_o21ai_1
X_2260_ net919 controller.counter2.counter_0\[1\] controller.counter2.counter_0\[0\]
+ _0406_ VPWR VGND sg13g2_nor3_1
XFILLER_33_386 VPWR VGND sg13g2_fill_2
X_1975_ net628 VPWR _1314_ VGND controller.inst_mem.mem_data\[85\] net555 sg13g2_o21ai_1
X_2458_ _0601_ net463 _0545_ VPWR VGND sg13g2_nand2b_1
X_2527_ _0651_ net954 _0657_ VPWR VGND sg13g2_xor2_1
Xhold16 _0013_ VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold27 _0142_ VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold38 _0138_ VPWR VGND net365 sg13g2_dlygate4sd3_1
X_2389_ VPWR VGND controller.inst_mem.mem_data\[150\] net517 net520 controller.inst_mem.mem_data\[102\]
+ _0532_ net495 sg13g2_a221oi_1
Xhold49 controller.extended_state\[0\] VPWR VGND net376 sg13g2_dlygate4sd3_1
X_3133__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_47_401 VPWR VGND sg13g2_decap_8
XFILLER_47_478 VPWR VGND sg13g2_decap_8
X_1691_ VPWR _1042_ net409 VGND sg13g2_inv_1
XFILLER_30_323 VPWR VGND sg13g2_fill_1
X_1760_ VPWR _1111_ net430 VGND sg13g2_inv_1
X_2312_ _0448_ _0457_ _0458_ VPWR VGND sg13g2_nor2b_1
X_2174_ VGND VPWR _1113_ net546 _0103_ _0362_ sg13g2_a21oi_1
X_2243_ net651 VPWR _0397_ VGND controller.inst_mem.extended_word\[19\] net602 sg13g2_o21ai_1
Xoutput17 net17 uo_out[2] VPWR VGND sg13g2_buf_1
X_1889_ _1240_ _1237_ _1239_ VPWR VGND sg13g2_nand2_1
X_1958_ _1304_ _1258_ controller.alu_buffer.buffer\[5\] _1257_ net536 VPWR VGND sg13g2_a22oi_1
XFILLER_44_415 VPWR VGND sg13g2_decap_8
X_3142__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_43_492 VPWR VGND sg13g2_decap_8
X_2861_ net658 VPWR _0922_ VGND net820 net614 sg13g2_o21ai_1
X_2930_ VGND VPWR _1004_ net587 _0265_ _0956_ sg13g2_a21oi_1
Xhold349 controller.counter2.counter_0\[8\] VPWR VGND net896 sg13g2_dlygate4sd3_1
X_2792_ _1277_ net942 _0880_ VPWR VGND sg13g2_xor2_1
Xhold305 controller.inst_mem.mem_data\[49\] VPWR VGND net852 sg13g2_dlygate4sd3_1
Xhold338 controller.extended_cond.opcode\[2\] VPWR VGND net885 sg13g2_dlygate4sd3_1
Xhold316 controller.inst_mem.mem_data\[182\] VPWR VGND net863 sg13g2_dlygate4sd3_1
X_1812_ VPWR _1163_ net384 VGND sg13g2_inv_1
X_1743_ VPWR _1094_ net842 VGND sg13g2_inv_1
X_1674_ VPWR _1025_ net748 VGND sg13g2_inv_1
Xhold327 controller.inst_mem.mem_data\[78\] VPWR VGND net874 sg13g2_dlygate4sd3_1
XFILLER_30_0 VPWR VGND sg13g2_fill_1
X_2226_ VGND VPWR _1087_ net575 _0129_ _0388_ sg13g2_a21oi_1
X_3086__241 VPWR VGND net241 sg13g2_tiehi
X_2157_ net649 VPWR _0354_ VGND controller.inst_mem.mem_data\[176\] net594 sg13g2_o21ai_1
X_2088_ VGND VPWR _1156_ net590 _0060_ _0319_ sg13g2_a21oi_1
XFILLER_34_492 VPWR VGND sg13g2_decap_8
XFILLER_21_153 VPWR VGND sg13g2_fill_2
XFILLER_44_201 VPWR VGND sg13g2_fill_2
XFILLER_40_462 VPWR VGND sg13g2_decap_8
XFILLER_12_131 VPWR VGND sg13g2_fill_1
XFILLER_17_459 VPWR VGND sg13g2_fill_1
X_2998__128 VPWR VGND net128 sg13g2_tiehi
X_3060_ net293 VGND VPWR _0083_ controller.inst_mem.mem_data\[164\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_2011_ net649 VPWR _1332_ VGND controller.inst_mem.mem_data\[103\] net595 sg13g2_o21ai_1
X_2844_ VGND VPWR _1047_ net577 _0222_ _0913_ sg13g2_a21oi_1
X_2913_ net657 VPWR _0948_ VGND controller.inst_mem.mem_data\[49\] net610 sg13g2_o21ai_1
X_3036__52 VPWR VGND net52 sg13g2_tiehi
Xhold168 controller.const_data\[6\] VPWR VGND net715 sg13g2_dlygate4sd3_1
Xhold124 controller.const_data\[0\] VPWR VGND net671 sg13g2_dlygate4sd3_1
X_2775_ VGND VPWR net476 _0865_ _0200_ _0866_ sg13g2_a21oi_1
Xhold113 controller.const_data\[29\] VPWR VGND net440 sg13g2_dlygate4sd3_1
X_1726_ VPWR _1077_ net392 VGND sg13g2_inv_1
Xhold146 controller.inst_mem.mem_data\[44\] VPWR VGND net693 sg13g2_dlygate4sd3_1
Xhold135 controller.inst_mem.mem_data\[193\] VPWR VGND net682 sg13g2_dlygate4sd3_1
Xfanout615 net616 net615 VPWR VGND sg13g2_buf_8
Xhold157 _0075_ VPWR VGND net704 sg13g2_dlygate4sd3_1
Xhold102 _0054_ VPWR VGND net429 sg13g2_dlygate4sd3_1
X_1657_ VPWR _1008_ net786 VGND sg13g2_inv_1
Xhold179 controller.inst_mem.mem_data\[54\] VPWR VGND net726 sg13g2_dlygate4sd3_1
Xfanout604 net605 net604 VPWR VGND sg13g2_buf_2
X_3189_ net196 VGND VPWR _0212_ controller.const_data\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_1
Xfanout637 net663 net637 VPWR VGND sg13g2_buf_8
Xfanout659 net663 net659 VPWR VGND sg13g2_buf_8
X_3258_ net147 VGND VPWR _0281_ controller.inst_mem.mem_data\[73\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_2209_ net645 VPWR _0380_ VGND net842 net583 sg13g2_o21ai_1
Xfanout648 net650 net648 VPWR VGND sg13g2_buf_8
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_8
X_2491_ _0628_ net457 net12 net472 net961 VPWR VGND sg13g2_a22oi_1
X_2560_ VGND VPWR _0682_ _0683_ _0167_ _0684_ sg13g2_a21oi_1
X_3112_ net189 VGND VPWR _0135_ controller.extended_then_action\[4\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_3043_ net327 VGND VPWR _0066_ controller.inst_mem.mem_data\[147\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_2827_ net636 VPWR _0905_ VGND net715 net569 sg13g2_o21ai_1
X_2758_ VGND VPWR net718 net453 _0853_ _0852_ sg13g2_a21oi_1
X_3170__272 VPWR VGND net272 sg13g2_tiehi
X_2689_ VPWR VGND net13 net446 _0774_ net715 _0799_ net479 sg13g2_a221oi_1
X_1709_ VPWR _1060_ net671 VGND sg13g2_inv_1
Xfanout445 _0773_ net445 VPWR VGND sg13g2_buf_8
Xfanout456 net457 net456 VPWR VGND sg13g2_buf_8
X_3129__141 VPWR VGND net141 sg13g2_tiehi
Xfanout478 _0748_ net478 VPWR VGND sg13g2_buf_2
Xfanout467 net469 net467 VPWR VGND sg13g2_buf_8
Xfanout489 _0438_ net489 VPWR VGND sg13g2_buf_2
XFILLER_10_421 VPWR VGND sg13g2_fill_2
XFILLER_38_81 VPWR VGND sg13g2_fill_2
X_2612_ _0727_ VPWR _0728_ VGND controller.inst_mem.mem_data\[45\] net492 sg13g2_o21ai_1
X_1991_ net655 VPWR _1322_ VGND net342 net607 sg13g2_o21ai_1
Xclkload11 VPWR clkload11/Y clknet_leaf_22_clk VGND sg13g2_inv_1
X_2474_ _0614_ _0612_ _0613_ VPWR VGND sg13g2_nand2_1
X_2543_ controller.alu_buffer.buffer\[16\] _1294_ _0670_ VPWR VGND sg13g2_and2_1
X_3026_ net72 VGND VPWR net341 controller.inst_mem.mem_data\[130\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
Xclkload5 clkload5/Y clknet_leaf_12_clk VPWR VGND sg13g2_inv_2
X_3184__216 VPWR VGND net216 sg13g2_tiehi
X_2190_ VGND VPWR _1105_ net617 _0111_ _0370_ sg13g2_a21oi_1
X_1974_ VGND VPWR _1213_ net559 _0003_ _1313_ sg13g2_a21oi_1
X_3045__323 VPWR VGND net323 sg13g2_tiehi
Xhold17 controller.const_data\[19\] VPWR VGND net344 sg13g2_dlygate4sd3_1
X_2457_ _0599_ _0585_ _0563_ _0600_ VPWR VGND sg13g2_a21o_1
X_2526_ controller.alu_buffer.buffer\[13\] controller.alu_buffer.buffer\[12\] _1291_
+ _0656_ VPWR VGND sg13g2_nor3_1
Xhold39 controller.inst_mem.mem_data\[74\] VPWR VGND net366 sg13g2_dlygate4sd3_1
X_2388_ _0531_ net503 controller.inst_mem.mem_data\[198\] net507 controller.inst_mem.mem_data\[78\]
+ VPWR VGND sg13g2_a22oi_1
Xhold28 controller.inst_mem.mem_data\[138\] VPWR VGND net355 sg13g2_dlygate4sd3_1
X_3009_ net106 VGND VPWR _0032_ controller.inst_mem.mem_data\[113\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_3096__221 VPWR VGND net221 sg13g2_tiehi
XFILLER_3_247 VPWR VGND sg13g2_fill_2
XFILLER_47_457 VPWR VGND sg13g2_decap_8
XFILLER_19_115 VPWR VGND sg13g2_fill_1
X_1690_ VPWR _1041_ net344 VGND sg13g2_inv_1
XFILLER_30_368 VPWR VGND sg13g2_fill_1
X_2242_ VGND VPWR _1079_ net615 _0137_ _0396_ sg13g2_a21oi_1
X_2311_ _0455_ _0450_ _0456_ _0457_ VPWR VGND sg13g2_a21o_2
XFILLER_46_490 VPWR VGND sg13g2_decap_8
XFILLER_38_479 VPWR VGND sg13g2_decap_8
X_2173_ net627 VPWR _0362_ VGND controller.inst_mem.mem_data\[184\] net546 sg13g2_o21ai_1
XFILLER_21_302 VPWR VGND sg13g2_fill_2
X_1957_ _1303_ controller.alu_buffer.buffer\[21\] _1260_ VPWR VGND sg13g2_nand2_1
X_2509_ _0642_ _1290_ _0641_ VPWR VGND sg13g2_nand2_1
Xoutput18 net18 uo_out[3] VPWR VGND sg13g2_buf_1
X_1888_ VPWR VGND controller.inst_mem.mem_data\[136\] net514 net519 controller.inst_mem.mem_data\[112\]
+ _1239_ net498 sg13g2_a221oi_1
Xclkbuf_leaf_36_clk clknet_3_1__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_12_324 VPWR VGND sg13g2_fill_2
XFILLER_47_276 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_27_clk clknet_3_5__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_43_471 VPWR VGND sg13g2_decap_8
X_2860_ VGND VPWR _1039_ net613 _0230_ _0921_ sg13g2_a21oi_1
X_2791_ VGND VPWR net478 _0878_ _0203_ _0879_ sg13g2_a21oi_1
X_1811_ VPWR _1162_ net428 VGND sg13g2_inv_1
Xhold339 controller.counter2.counter_0\[9\] VPWR VGND net886 sg13g2_dlygate4sd3_1
Xhold306 controller.inst_mem.mem_data\[43\] VPWR VGND net853 sg13g2_dlygate4sd3_1
Xhold328 controller.inst_mem.mem_data\[156\] VPWR VGND net875 sg13g2_dlygate4sd3_1
X_1673_ _1024_ net876 VPWR VGND sg13g2_inv_2
Xhold317 controller.inst_mem.mem_data\[61\] VPWR VGND net864 sg13g2_dlygate4sd3_1
X_1742_ VPWR _1093_ net729 VGND sg13g2_inv_1
X_2225_ net639 VPWR _0388_ VGND controller.extended_cond.opcode\[1\] net575 sg13g2_o21ai_1
XFILLER_23_0 VPWR VGND sg13g2_fill_2
XFILLER_34_471 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_3_7__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_2156_ VGND VPWR _1122_ net595 _0094_ _0353_ sg13g2_a21oi_1
X_2087_ net646 VPWR _0319_ VGND net330 net590 sg13g2_o21ai_1
X_2989_ net146 VGND VPWR _0012_ controller.inst_mem.mem_data\[93\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
XFILLER_40_441 VPWR VGND sg13g2_decap_8
X_3102__209 VPWR VGND net209 sg13g2_tiehi
X_2010_ VGND VPWR _1195_ net595 _0021_ _1331_ sg13g2_a21oi_1
X_2912_ VGND VPWR _1013_ net607 _0256_ _0947_ sg13g2_a21oi_1
X_2843_ net640 VPWR _0913_ VGND net694 net577 sg13g2_o21ai_1
X_2774_ net543 VPWR _0866_ VGND net921 net476 sg13g2_o21ai_1
X_1725_ VPWR _1076_ net403 VGND sg13g2_inv_1
XFILLER_31_463 VPWR VGND sg13g2_fill_2
X_3003__118 VPWR VGND net118 sg13g2_tiehi
Xhold147 controller.const_data\[14\] VPWR VGND net694 sg13g2_dlygate4sd3_1
Xhold169 _0215_ VPWR VGND net716 sg13g2_dlygate4sd3_1
Xhold125 _0209_ VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold114 _0238_ VPWR VGND net441 sg13g2_dlygate4sd3_1
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_7_clk clknet_3_2__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xfanout616 net622 net616 VPWR VGND sg13g2_buf_8
Xhold158 controller.inst_mem.mem_data\[81\] VPWR VGND net705 sg13g2_dlygate4sd3_1
Xfanout649 net650 net649 VPWR VGND sg13g2_buf_8
Xfanout627 net635 net627 VPWR VGND sg13g2_buf_8
X_1656_ VPWR _1007_ net812 VGND sg13g2_inv_1
Xfanout605 net624 net605 VPWR VGND sg13g2_buf_8
Xhold136 controller.inst_mem.extended_word\[21\] VPWR VGND net683 sg13g2_dlygate4sd3_1
Xhold103 controller.inst_mem.mem_data\[185\] VPWR VGND net430 sg13g2_dlygate4sd3_1
X_3188_ net200 VGND VPWR net833 controller.const_data\[3\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3257_ net190 VGND VPWR net670 controller.inst_mem.mem_data\[72\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
XFILLER_26_246 VPWR VGND sg13g2_fill_1
X_2139_ net656 VPWR _0345_ VGND net350 net608 sg13g2_o21ai_1
X_2208_ VGND VPWR _1096_ net587 _0120_ _0379_ sg13g2_a21oi_1
XFILLER_5_139 VPWR VGND sg13g2_fill_1
X_2490_ VPWR VGND net469 net464 _0626_ net527 _0627_ net483 sg13g2_a221oi_1
XFILLER_48_393 VPWR VGND sg13g2_decap_8
X_3111_ net191 VGND VPWR net686 controller.extended_then_action\[3\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_3042_ net40 VGND VPWR net680 controller.inst_mem.mem_data\[146\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_3159__316 VPWR VGND net316 sg13g2_tiehi
X_1708_ VPWR _1059_ net695 VGND sg13g2_inv_1
X_2757_ VGND VPWR _1271_ _0851_ _0852_ net452 sg13g2_a21oi_1
X_2688_ net448 VPWR _0798_ VGND _0410_ _0797_ sg13g2_o21ai_1
X_2826_ VGND VPWR _1056_ net569 _0213_ _0904_ sg13g2_a21oi_1
X_3055__303 VPWR VGND net303 sg13g2_tiehi
Xfanout446 net447 net446 VPWR VGND sg13g2_buf_8
Xfanout479 net480 net479 VPWR VGND sg13g2_buf_8
Xfanout468 net469 net468 VPWR VGND sg13g2_buf_8
Xfanout457 _0607_ net457 VPWR VGND sg13g2_buf_8
X_1639_ VPWR _0990_ net803 VGND sg13g2_inv_1
X_3263__45 VPWR VGND net45 sg13g2_tiehi
X_3136__113 VPWR VGND net113 sg13g2_tiehi
X_1990_ VGND VPWR _1205_ net567 _0011_ _1321_ sg13g2_a21oi_1
X_2611_ _0724_ _0725_ _0723_ _0727_ VPWR VGND _0726_ sg13g2_nand4_1
X_2542_ controller.alu_buffer.buffer\[16\] _1294_ _0669_ VPWR VGND sg13g2_nor2_1
X_2473_ net529 VPWR _0613_ VGND net530 net984 sg13g2_o21ai_1
X_3230__178 VPWR VGND net178 sg13g2_tiehi
X_3025_ net74 VGND VPWR _0048_ controller.inst_mem.mem_data\[129\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_2987__150 VPWR VGND net150 sg13g2_tiehi
X_3198__151 VPWR VGND net151 sg13g2_tiehi
Xclkload6 VPWR clkload6/Y clknet_leaf_13_clk VGND sg13g2_inv_1
X_2809_ VGND VPWR net474 _0893_ _0206_ _0894_ sg13g2_a21oi_1
X_1973_ net630 VPWR _1313_ VGND net724 net559 sg13g2_o21ai_1
X_2525_ VPWR VGND net950 net462 net482 controller.alu_buffer.buffer\[12\] _0655_ net471
+ sg13g2_a221oi_1
Xhold18 _0228_ VPWR VGND net345 sg13g2_dlygate4sd3_1
X_2456_ VPWR VGND _0597_ _0598_ net463 net468 _0599_ _0587_ sg13g2_a221oi_1
X_2387_ _0530_ net499 controller.inst_mem.mem_data\[126\] net511 controller.inst_mem.mem_data\[174\]
+ VPWR VGND sg13g2_a22oi_1
Xhold29 _0058_ VPWR VGND net356 sg13g2_dlygate4sd3_1
XFILLER_28_149 VPWR VGND sg13g2_fill_1
X_3008_ net108 VGND VPWR net731 controller.inst_mem.mem_data\[112\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_47_436 VPWR VGND sg13g2_decap_8
X_2172_ VGND VPWR _1114_ net546 _0102_ _0361_ sg13g2_a21oi_1
X_3145__77 VPWR VGND net77 sg13g2_tiehi
X_2310_ controller.inst_mem.mem_data\[43\] net493 _0456_ VPWR VGND sg13g2_nor2_1
X_2241_ net661 VPWR _0396_ VGND net364 net615 sg13g2_o21ai_1
XFILLER_38_458 VPWR VGND sg13g2_decap_8
XFILLER_33_163 VPWR VGND sg13g2_fill_2
XFILLER_18_171 VPWR VGND sg13g2_fill_2
XFILLER_18_182 VPWR VGND sg13g2_fill_1
X_1956_ net19 _1301_ _1302_ VPWR VGND sg13g2_nand2_2
X_1887_ _1238_ net494 controller.inst_mem.mem_data\[88\] net502 controller.inst_mem.mem_data\[184\]
+ VPWR VGND sg13g2_a22oi_1
X_2508_ controller.alu_buffer.buffer\[10\] VPWR _0641_ VGND controller.alu_buffer.buffer\[9\]
+ _1288_ sg13g2_o21ai_1
Xoutput19 net19 uo_out[4] VPWR VGND sg13g2_buf_1
X_2439_ _0582_ _0573_ _0580_ VPWR VGND sg13g2_nand2_2
X_3063__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_12_369 VPWR VGND sg13g2_fill_1
XFILLER_20_380 VPWR VGND sg13g2_fill_2
XFILLER_43_450 VPWR VGND sg13g2_decap_8
X_2790_ net543 VPWR _0879_ VGND net883 net478 sg13g2_o21ai_1
X_1810_ VPWR _1161_ net668 VGND sg13g2_inv_1
X_3109__195 VPWR VGND net195 sg13g2_tiehi
X_1741_ VPWR _1092_ net334 VGND sg13g2_inv_1
X_1672_ VPWR _1023_ net869 VGND sg13g2_inv_1
Xhold318 controller.inst_mem.mem_data\[102\] VPWR VGND net865 sg13g2_dlygate4sd3_1
Xhold329 controller.inst_mem.mem_data\[36\] VPWR VGND net876 sg13g2_dlygate4sd3_1
Xhold307 controller.extended_jump_target\[1\] VPWR VGND net854 sg13g2_dlygate4sd3_1
XFILLER_38_244 VPWR VGND sg13g2_fill_2
X_2155_ net649 VPWR _0353_ VGND net699 net597 sg13g2_o21ai_1
X_2224_ VGND VPWR _1088_ net554 _0128_ _0387_ sg13g2_a21oi_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
X_2086_ VGND VPWR _1157_ net565 _0059_ _0318_ sg13g2_a21oi_1
X_1939_ controller.alu_buffer.buffer\[7\] net527 _1286_ VPWR VGND sg13g2_nor2_1
X_2988_ net148 VGND VPWR net443 controller.inst_mem.mem_data\[92\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_3173__260 VPWR VGND net260 sg13g2_tiehi
XFILLER_40_497 VPWR VGND sg13g2_decap_8
X_3221__250 VPWR VGND net250 sg13g2_tiehi
XFILLER_8_159 VPWR VGND sg13g2_fill_1
X_2911_ net657 VPWR _0947_ VGND net407 net609 sg13g2_o21ai_1
X_2842_ VGND VPWR _1048_ net577 _0221_ _0912_ sg13g2_a21oi_1
X_2773_ VGND VPWR net811 net452 _0865_ _0864_ sg13g2_a21oi_1
XFILLER_31_486 VPWR VGND sg13g2_decap_8
X_1724_ VPWR _1075_ net683 VGND sg13g2_inv_1
Xhold115 controller.inst_mem.mem_data\[91\] VPWR VGND net442 sg13g2_dlygate4sd3_1
Xhold104 _0105_ VPWR VGND net431 sg13g2_dlygate4sd3_1
Xhold126 controller.inst_mem.mem_data\[116\] VPWR VGND net673 sg13g2_dlygate4sd3_1
Xhold148 controller.const_data\[1\] VPWR VGND net695 sg13g2_dlygate4sd3_1
X_3256_ net222 VGND VPWR _0279_ controller.inst_mem.mem_data\[71\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
Xfanout639 net641 net639 VPWR VGND sg13g2_buf_2
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_8
Xfanout617 net622 net617 VPWR VGND sg13g2_buf_8
Xhold159 controller.inst_mem.mem_data\[179\] VPWR VGND net706 sg13g2_dlygate4sd3_1
Xfanout628 net629 net628 VPWR VGND sg13g2_buf_8
X_1655_ VPWR _1006_ net726 VGND sg13g2_inv_1
Xhold137 controller.inst_mem.mem_data\[92\] VPWR VGND net684 sg13g2_dlygate4sd3_1
X_3187_ net204 VGND VPWR net696 controller.const_data\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2069_ net630 VPWR _0310_ VGND net692 net560 sg13g2_o21ai_1
X_2207_ net644 VPWR _0379_ VGND controller.extended_jump_target\[1\] net587 sg13g2_o21ai_1
X_2138_ VGND VPWR _1131_ net590 _0085_ _0344_ sg13g2_a21oi_1
XFILLER_41_217 VPWR VGND sg13g2_fill_1
X_2997__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_1_368 VPWR VGND sg13g2_fill_1
XFILLER_27_73 VPWR VGND sg13g2_fill_1
XFILLER_9_413 VPWR VGND sg13g2_fill_2
X_3187__204 VPWR VGND net204 sg13g2_tiehi
X_3110_ net193 VGND VPWR _0133_ controller.extended_then_action\[2\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
XFILLER_48_372 VPWR VGND sg13g2_decap_8
X_3041_ net42 VGND VPWR net333 controller.inst_mem.mem_data\[145\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_2825_ net636 VPWR _0904_ VGND controller.const_data\[5\] net569 sg13g2_o21ai_1
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_2756_ net910 VPWR _0851_ VGND net903 _1270_ sg13g2_o21ai_1
X_2687_ _0409_ net894 _0797_ VPWR VGND sg13g2_nor2b_1
X_1707_ VPWR _1058_ net832 VGND sg13g2_inv_1
X_1638_ VPWR _0989_ net669 VGND sg13g2_inv_1
Xfanout447 _0772_ net447 VPWR VGND sg13g2_buf_8
Xfanout469 _0586_ net469 VPWR VGND sg13g2_buf_2
Xfanout458 net459 net458 VPWR VGND sg13g2_buf_8
X_3239_ net326 VGND VPWR _0262_ controller.inst_mem.mem_data\[54\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_10_445 VPWR VGND sg13g2_fill_2
XFILLER_22_294 VPWR VGND sg13g2_fill_2
XFILLER_45_364 VPWR VGND sg13g2_fill_2
X_2472_ net529 net530 net984 _0612_ VPWR VGND sg13g2_or3_1
X_2541_ controller.alu_buffer.buffer\[8\] _0562_ _0668_ VPWR VGND sg13g2_nor2_1
X_2610_ VGND VPWR controller.inst_mem.mem_data\[189\] net502 _0726_ net515 sg13g2_a21oi_1
XFILLER_36_397 VPWR VGND sg13g2_fill_2
X_3024_ net76 VGND VPWR _0047_ controller.inst_mem.mem_data\[128\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_2808_ net544 VPWR _0894_ VGND net904 net474 sg13g2_o21ai_1
Xclkload7 clkload7/Y clknet_leaf_31_clk VPWR VGND sg13g2_inv_2
X_2739_ VGND VPWR net475 _0836_ _0193_ _0837_ sg13g2_a21oi_1
XFILLER_30_507 VPWR VGND sg13g2_fill_1
XFILLER_24_85 VPWR VGND sg13g2_fill_1
X_3073__267 VPWR VGND net267 sg13g2_tiehi
X_1972_ VGND VPWR _1214_ net581 _0002_ _1312_ sg13g2_a21oi_1
XFILLER_46_0 VPWR VGND sg13g2_fill_1
X_2455_ VGND VPWR _1065_ _0561_ _0598_ net485 sg13g2_a21oi_1
X_2524_ VGND VPWR _0650_ _0653_ _0161_ _0654_ sg13g2_a21oi_1
X_3119__175 VPWR VGND net175 sg13g2_tiehi
Xhold19 controller.inst_mem.mem_data\[73\] VPWR VGND net346 sg13g2_dlygate4sd3_1
X_2386_ _0529_ controller.inst_mem.extended_word\[22\] net524 VPWR VGND sg13g2_nand2_1
X_3007_ net110 VGND VPWR _0030_ controller.inst_mem.mem_data\[111\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_47_415 VPWR VGND sg13g2_decap_8
X_2240_ VGND VPWR _1080_ net616 _0136_ _0395_ sg13g2_a21oi_1
X_2171_ net627 VPWR _0361_ VGND net378 net547 sg13g2_o21ai_1
X_1955_ _1302_ _1299_ _1257_ _1258_ net528 VPWR VGND sg13g2_a22oi_1
X_1886_ _1237_ controller.inst_mem.mem_data\[64\] net506 VPWR VGND sg13g2_nand2_1
XFILLER_21_359 VPWR VGND sg13g2_fill_1
X_2507_ VPWR VGND _0640_ _0503_ _0638_ _1065_ _0158_ net463 sg13g2_a221oi_1
X_2438_ _0573_ _0580_ _0581_ VPWR VGND sg13g2_and2_1
XFILLER_44_429 VPWR VGND sg13g2_decap_8
X_2369_ net486 _0511_ _0514_ VPWR VGND sg13g2_nor2_1
XFILLER_24_186 VPWR VGND sg13g2_fill_1
XFILLER_47_278 VPWR VGND sg13g2_fill_1
X_1740_ VPWR _1091_ net710 VGND sg13g2_inv_1
Xhold308 controller.inst_mem.mem_data\[109\] VPWR VGND net855 sg13g2_dlygate4sd3_1
X_1671_ VPWR _1022_ net877 VGND sg13g2_inv_1
Xhold319 _0022_ VPWR VGND net866 sg13g2_dlygate4sd3_1
X_2154_ VGND VPWR _1123_ net596 _0093_ _0352_ sg13g2_a21oi_1
X_2223_ net632 VPWR _0387_ VGND controller.extended_cond.opcode\[0\] net554 sg13g2_o21ai_1
X_2085_ net633 VPWR _0318_ VGND controller.inst_mem.mem_data\[140\] net565 sg13g2_o21ai_1
X_2987_ net150 VGND VPWR net424 controller.inst_mem.mem_data\[91\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_1938_ _1285_ _1283_ _1284_ VPWR VGND sg13g2_nand2_2
X_3211__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_1_506 VPWR VGND sg13g2_fill_2
X_1869_ _1068_ _1216_ _1220_ VPWR VGND sg13g2_and2_1
X_3180__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_40_476 VPWR VGND sg13g2_decap_8
X_3139__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_35_215 VPWR VGND sg13g2_fill_1
X_2841_ net640 VPWR _0912_ VGND controller.const_data\[13\] net577 sg13g2_o21ai_1
X_2910_ VGND VPWR _1014_ net606 _0255_ _0946_ sg13g2_a21oi_1
Xhold149 _0210_ VPWR VGND net696 sg13g2_dlygate4sd3_1
X_2772_ net452 _0863_ _0864_ VPWR VGND sg13g2_nor2_1
Xhold138 controller.extended_then_action\[2\] VPWR VGND net685 sg13g2_dlygate4sd3_1
X_1654_ VPWR _1005_ net872 VGND sg13g2_inv_1
X_1723_ VPWR _1074_ net353 VGND sg13g2_inv_1
Xhold116 _0011_ VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold105 controller.inst_mem.mem_data\[51\] VPWR VGND net432 sg13g2_dlygate4sd3_1
Xhold127 _0036_ VPWR VGND net674 sg13g2_dlygate4sd3_1
Xfanout618 net622 net618 VPWR VGND sg13g2_buf_1
Xfanout607 net623 net607 VPWR VGND sg13g2_buf_8
X_3255_ net254 VGND VPWR _0278_ controller.inst_mem.mem_data\[70\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
Xfanout629 net631 net629 VPWR VGND sg13g2_buf_8
X_2206_ VGND VPWR _1097_ net593 _0119_ _0378_ sg13g2_a21oi_1
X_3186_ net208 VGND VPWR net672 controller.const_data\[1\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_2137_ net655 VPWR _0344_ VGND controller.inst_mem.mem_data\[166\] net607 sg13g2_o21ai_1
X_2068_ VGND VPWR _1166_ net584 _0050_ _0309_ sg13g2_a21oi_1
X_3101__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_22_498 VPWR VGND sg13g2_fill_1
XFILLER_1_358 VPWR VGND sg13g2_fill_2
X_3018__88 VPWR VGND net88 sg13g2_tiehi
X_3002__120 VPWR VGND net120 sg13g2_tiehi
X_3033__58 VPWR VGND net58 sg13g2_tiehi
X_3083__247 VPWR VGND net247 sg13g2_tiehi
X_3040_ net44 VGND VPWR _0063_ controller.inst_mem.mem_data\[144\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_2824_ VGND VPWR _1057_ net569 _0212_ _0903_ sg13g2_a21oi_1
X_2755_ VGND VPWR net476 _0849_ _0196_ _0850_ sg13g2_a21oi_1
X_2686_ VGND VPWR _0794_ _0795_ _0181_ _0796_ sg13g2_a21oi_1
X_1706_ VPWR _1057_ net838 VGND sg13g2_inv_1
X_1637_ VPWR _0988_ net734 VGND sg13g2_inv_1
Xfanout448 net449 net448 VPWR VGND sg13g2_buf_8
X_3169_ net276 VGND VPWR _0192_ controller.counter2.counter_1\[0\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
Xfanout459 _0596_ net459 VPWR VGND sg13g2_buf_8
X_3238_ net59 VGND VPWR net787 controller.inst_mem.mem_data\[53\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_42_505 VPWR VGND sg13g2_fill_2
XFILLER_6_428 VPWR VGND sg13g2_fill_1
XFILLER_10_413 VPWR VGND sg13g2_fill_2
X_2471_ VPWR VGND net977 net463 net483 net530 _0611_ net472 sg13g2_a221oi_1
X_2540_ VPWR VGND _0667_ _0503_ _0665_ _1064_ _0164_ net461 sg13g2_a221oi_1
X_3023_ net78 VGND VPWR net667 controller.inst_mem.mem_data\[127\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_2738_ net544 VPWR _0837_ VGND net915 net475 sg13g2_o21ai_1
X_2807_ VGND VPWR net689 net450 _0893_ _0892_ sg13g2_a21oi_1
Xclkload8 VPWR clkload8/Y clknet_leaf_32_clk VGND sg13g2_inv_1
X_2669_ VPWR VGND net9 net446 _0774_ net832 _0783_ net479 sg13g2_a221oi_1
XFILLER_27_332 VPWR VGND sg13g2_fill_1
XFILLER_27_398 VPWR VGND sg13g2_fill_1
XFILLER_40_74 VPWR VGND sg13g2_fill_1
XFILLER_6_0 VPWR VGND sg13g2_fill_1
XFILLER_45_162 VPWR VGND sg13g2_fill_1
X_1971_ net642 VPWR _1312_ VGND controller.inst_mem.mem_data\[83\] net581 sg13g2_o21ai_1
X_2454_ net485 _0594_ _0597_ VPWR VGND sg13g2_and2_1
X_3148__65 VPWR VGND net65 sg13g2_tiehi
X_2523_ net538 VPWR _0654_ VGND net969 net459 sg13g2_o21ai_1
X_2385_ _1080_ net490 net489 _0528_ VPWR VGND sg13g2_or3_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_3006_ net112 VGND VPWR _0029_ controller.inst_mem.mem_data\[110\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_42_121 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_39_clk clknet_3_0__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
X_2170_ VGND VPWR _1115_ net548 _0101_ _0360_ sg13g2_a21oi_1
X_1954_ _1301_ controller.alu_buffer.buffer\[20\] _1260_ VPWR VGND sg13g2_nand2_1
X_1885_ VPWR _1236_ _1235_ VGND sg13g2_inv_1
X_2506_ _0640_ _0639_ net468 _0607_ controller.alu_buffer.buffer\[1\] VPWR VGND sg13g2_a22oi_1
X_2437_ VGND VPWR _0475_ _0579_ _0580_ _0485_ sg13g2_a21oi_1
X_2368_ _0505_ net488 _0512_ _0513_ VPWR VGND sg13g2_a21o_1
XFILLER_44_408 VPWR VGND sg13g2_decap_8
XFILLER_37_482 VPWR VGND sg13g2_decap_8
X_2299_ VPWR VGND controller.inst_mem.mem_data\[114\] _0443_ net498 controller.inst_mem.mem_data\[66\]
+ _0445_ net509 sg13g2_a221oi_1
X_3254__286 VPWR VGND net286 sg13g2_tiehi
XFILLER_43_485 VPWR VGND sg13g2_decap_8
XFILLER_30_135 VPWR VGND sg13g2_fill_2
X_1670_ VPWR _1021_ net799 VGND sg13g2_inv_1
Xhold309 controller.inst_mem.mem_data\[41\] VPWR VGND net856 sg13g2_dlygate4sd3_1
X_2222_ VGND VPWR _1089_ net551 _0127_ _0386_ sg13g2_a21oi_1
X_3012__100 VPWR VGND net100 sg13g2_tiehi
X_3141__93 VPWR VGND net93 sg13g2_tiehi
X_2153_ net650 VPWR _0352_ VGND net738 net597 sg13g2_o21ai_1
X_2084_ VGND VPWR _1158_ net566 _0058_ _0317_ sg13g2_a21oi_1
X_1937_ controller.alu_buffer.buffer\[5\] net528 _1284_ VPWR VGND sg13g2_nor2_1
XFILLER_34_485 VPWR VGND sg13g2_decap_8
X_2986_ net152 VGND VPWR _0009_ controller.inst_mem.mem_data\[90\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_1868_ _1219_ controller.inst_mem.mem_data\[159\] net510 VPWR VGND sg13g2_nand2_1
X_3093__227 VPWR VGND net227 sg13g2_tiehi
X_1799_ VPWR _1150_ net806 VGND sg13g2_inv_1
XFILLER_12_102 VPWR VGND sg13g2_fill_1
XFILLER_40_455 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_fill_2
XFILLER_16_430 VPWR VGND sg13g2_fill_1
X_2840_ VGND VPWR _1049_ net577 _0220_ _0911_ sg13g2_a21oi_1
XFILLER_43_260 VPWR VGND sg13g2_fill_1
X_2771_ _1273_ net921 _0863_ VPWR VGND sg13g2_xor2_1
Xhold117 controller.inst_mem.mem_data\[45\] VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold139 _0134_ VPWR VGND net686 sg13g2_dlygate4sd3_1
Xhold128 controller.inst_mem.mem_data\[68\] VPWR VGND net675 sg13g2_dlygate4sd3_1
X_1653_ VPWR _1004_ net804 VGND sg13g2_inv_1
X_1722_ VPWR _1073_ net783 VGND sg13g2_inv_1
Xhold106 _0260_ VPWR VGND net433 sg13g2_dlygate4sd3_1
X_3185_ net212 VGND VPWR _0208_ controller.const_data\[0\] clknet_leaf_13_clk sg13g2_dfrbpq_2
Xfanout619 net621 net619 VPWR VGND sg13g2_buf_8
Xfanout608 net611 net608 VPWR VGND sg13g2_buf_8
X_3254_ net286 VGND VPWR net676 controller.inst_mem.mem_data\[69\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_2205_ net648 VPWR _0378_ VGND controller.extended_jump_target\[0\] net593 sg13g2_o21ai_1
X_2067_ net642 VPWR _0309_ VGND controller.inst_mem.mem_data\[131\] net581 sg13g2_o21ai_1
X_2136_ VGND VPWR _1132_ net565 _0084_ _0343_ sg13g2_a21oi_1
X_2969_ net652 VPWR _0976_ VGND net826 net600 sg13g2_o21ai_1
X_3249__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_43_52 VPWR VGND sg13g2_fill_1
XFILLER_36_503 VPWR VGND sg13g2_decap_4
X_2823_ net636 VPWR _0903_ VGND net419 net569 sg13g2_o21ai_1
X_2754_ net544 VPWR _0850_ VGND net903 net476 sg13g2_o21ai_1
X_1705_ VPWR _1056_ net419 VGND sg13g2_inv_1
X_2685_ net540 VPWR _0796_ VGND net938 net444 sg13g2_o21ai_1
X_1636_ VPWR _0987_ net346 VGND sg13g2_inv_1
Xfanout449 _0770_ net449 VPWR VGND sg13g2_buf_8
X_3168_ net280 VGND VPWR _0191_ controller.counter2.counter_0\[15\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
XFILLER_39_396 VPWR VGND sg13g2_fill_2
X_2119_ net628 VPWR _0335_ VGND net867 net555 sg13g2_o21ai_1
X_3237_ net75 VGND VPWR net433 controller.inst_mem.mem_data\[52\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_3099_ net215 VGND VPWR _0122_ controller.inst_mem.extended_word\[3\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_3253__318 VPWR VGND net318 sg13g2_tiehi
XFILLER_10_469 VPWR VGND sg13g2_fill_2
XFILLER_38_63 VPWR VGND sg13g2_fill_2
XFILLER_45_311 VPWR VGND sg13g2_fill_1
XFILLER_9_278 VPWR VGND sg13g2_fill_1
X_2470_ VGND VPWR _0608_ _0609_ _0151_ _0610_ sg13g2_a21oi_1
XFILLER_36_322 VPWR VGND sg13g2_fill_2
X_3022_ net80 VGND VPWR net383 controller.inst_mem.mem_data\[126\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_2737_ VGND VPWR net410 net454 _0836_ _0835_ sg13g2_a21oi_1
X_2668_ net448 VPWR _0782_ VGND _0406_ _0781_ sg13g2_o21ai_1
X_2806_ net450 _0891_ _0892_ VPWR VGND sg13g2_nor2_1
Xclkload9 clknet_leaf_27_clk clkload9/X VPWR VGND sg13g2_buf_8
X_3020__84 VPWR VGND net84 sg13g2_tiehi
X_2599_ _0715_ net525 controller.inst_mem.extended_word\[19\] net511 controller.inst_mem.mem_data\[171\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_10_211 VPWR VGND sg13g2_fill_1
XFILLER_6_248 VPWR VGND sg13g2_fill_2
XFILLER_37_119 VPWR VGND sg13g2_fill_2
X_1970_ VGND VPWR _1215_ net586 _0001_ _1311_ sg13g2_a21oi_1
X_2522_ _0653_ _0652_ net467 net456 net528 VPWR VGND sg13g2_a22oi_1
X_2453_ _0596_ _0582_ VPWR VGND _0561_ sg13g2_nand2b_2
X_3052__309 VPWR VGND net309 sg13g2_tiehi
X_2384_ VGND VPWR _1068_ _0494_ _0148_ _0527_ sg13g2_a21oi_1
XFILLER_49_480 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
XFILLER_28_119 VPWR VGND sg13g2_fill_2
X_3005_ net114 VGND VPWR _0028_ controller.inst_mem.mem_data\[109\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_3_207 VPWR VGND sg13g2_fill_1
X_3154__47 VPWR VGND net47 sg13g2_tiehi
X_3183__220 VPWR VGND net220 sg13g2_tiehi
XFILLER_30_317 VPWR VGND sg13g2_fill_1
X_3162__304 VPWR VGND net304 sg13g2_tiehi
XFILLER_46_483 VPWR VGND sg13g2_decap_8
X_2984__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_18_130 VPWR VGND sg13g2_fill_1
X_1953_ _1296_ _1298_ _1300_ VPWR VGND controller.alu_buffer.buffer\[20\] sg13g2_nand3b_1
X_1884_ _1234_ VPWR _1235_ VGND controller.inst_mem.mem_data\[39\] net493 sg13g2_o21ai_1
XFILLER_21_317 VPWR VGND sg13g2_fill_1
X_2505_ _0639_ net963 _1288_ VPWR VGND sg13g2_xnor2_1
X_2436_ _0578_ VPWR _0579_ VGND controller.inst_mem.mem_data\[47\] net492 sg13g2_o21ai_1
XFILLER_29_406 VPWR VGND sg13g2_fill_1
X_2367_ net486 VPWR _0512_ VGND net854 net488 sg13g2_o21ai_1
X_2298_ controller.inst_mem.mem_data\[138\] net519 _0444_ VPWR VGND sg13g2_and2_1
XFILLER_37_461 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_fill_1
XFILLER_43_464 VPWR VGND sg13g2_decap_8
XFILLER_15_188 VPWR VGND sg13g2_fill_1
X_3205__95 VPWR VGND net95 sg13g2_tiehi
X_2152_ VGND VPWR _1124_ net600 _0092_ _0351_ sg13g2_a21oi_1
X_2221_ net626 VPWR _0386_ VGND net761 net551 sg13g2_o21ai_1
XFILLER_34_464 VPWR VGND sg13g2_decap_8
X_2083_ net633 VPWR _0317_ VGND controller.inst_mem.mem_data\[139\] net566 sg13g2_o21ai_1
X_1936_ controller.alu_buffer.buffer\[3\] net529 net530 _1283_ VGND VPWR net971 sg13g2_nor4_2
X_2985_ net154 VGND VPWR net371 controller.inst_mem.mem_data\[89\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_1867_ net536 net532 _1218_ VPWR VGND net533 sg13g2_nand3b_1
X_1798_ VPWR _1149_ net436 VGND sg13g2_inv_1
X_2419_ VGND VPWR _0562_ _0561_ net485 sg13g2_or2_1
XFILLER_40_434 VPWR VGND sg13g2_decap_8
XFILLER_25_431 VPWR VGND sg13g2_fill_1
X_2770_ VGND VPWR net476 _0861_ _0199_ _0862_ sg13g2_a21oi_1
XFILLER_31_412 VPWR VGND sg13g2_fill_2
X_1721_ VPWR _1072_ net376 VGND sg13g2_inv_1
Xfanout609 net610 net609 VPWR VGND sg13g2_buf_8
Xhold118 _0254_ VPWR VGND net665 sg13g2_dlygate4sd3_1
Xhold129 _0277_ VPWR VGND net676 sg13g2_dlygate4sd3_1
X_1652_ VPWR _1003_ net426 VGND sg13g2_inv_1
Xhold107 controller.inst_mem.mem_data\[50\] VPWR VGND net434 sg13g2_dlygate4sd3_1
XFILLER_39_501 VPWR VGND sg13g2_decap_8
X_3184_ net216 VGND VPWR _0207_ controller.counter2.counter_1\[15\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
X_2204_ VGND VPWR _1098_ net596 _0118_ _0377_ sg13g2_a21oi_1
XFILLER_14_0 VPWR VGND sg13g2_fill_1
X_2135_ net646 VPWR _0343_ VGND net359 net590 sg13g2_o21ai_1
X_3253_ net318 VGND VPWR _0276_ controller.inst_mem.mem_data\[68\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_2066_ VGND VPWR _1167_ net585 _0049_ _0308_ sg13g2_a21oi_1
X_2968_ VGND VPWR _0985_ net601 _0284_ _0975_ sg13g2_a21oi_1
X_2899_ net632 VPWR _0941_ VGND net740 net563 sg13g2_o21ai_1
X_1919_ _1268_ _1260_ controller.alu_buffer.buffer\[18\] _1258_ net529 VPWR VGND sg13g2_a22oi_1
XFILLER_48_386 VPWR VGND sg13g2_decap_8
XFILLER_16_272 VPWR VGND sg13g2_fill_1
XFILLER_23_209 VPWR VGND sg13g2_fill_1
X_2822_ VGND VPWR _1058_ net570 _0211_ _0902_ sg13g2_a21oi_1
X_1704_ VPWR _1055_ net774 VGND sg13g2_inv_1
X_2753_ VGND VPWR net736 net452 _0849_ _0848_ sg13g2_a21oi_1
X_2684_ VPWR VGND net12 net446 _0774_ net774 _0795_ net479 sg13g2_a221oi_1
X_3017__90 VPWR VGND net90 sg13g2_tiehi
X_3032__60 VPWR VGND net60 sg13g2_tiehi
X_1635_ VPWR _0986_ net366 VGND sg13g2_inv_1
XFILLER_42_507 VPWR VGND sg13g2_fill_1
X_3167_ net284 VGND VPWR _0190_ controller.counter2.counter_0\[14\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_2049_ net661 VPWR _0300_ VGND net362 net621 sg13g2_o21ai_1
X_2118_ VGND VPWR _1141_ net559 _0075_ _0334_ sg13g2_a21oi_1
X_3098_ net217 VGND VPWR _0121_ controller.extended_jump_target\[2\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
X_3236_ net91 VGND VPWR _0259_ controller.inst_mem.mem_data\[51\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_38_75 VPWR VGND sg13g2_fill_1
XFILLER_33_507 VPWR VGND sg13g2_fill_1
X_3158__320 VPWR VGND net320 sg13g2_tiehi
XFILLER_36_312 VPWR VGND sg13g2_fill_1
X_3009__106 VPWR VGND net106 sg13g2_tiehi
X_3021_ net82 VGND VPWR _0044_ controller.inst_mem.mem_data\[125\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_2805_ _0891_ net904 _0884_ VPWR VGND sg13g2_xnor2_1
X_2736_ net454 _0834_ _0835_ VPWR VGND sg13g2_nor2_1
X_3213__314 VPWR VGND net314 sg13g2_tiehi
X_2994__136 VPWR VGND net136 sg13g2_tiehi
X_2667_ _0405_ net919 _0781_ VPWR VGND sg13g2_nor2b_1
X_3059__295 VPWR VGND net295 sg13g2_tiehi
X_3219_ net266 VGND VPWR net721 controller.inst_mem.mem_data\[34\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2598_ net521 VPWR _0714_ VGND _1068_ controller.inst_mem.mem_data\[147\] sg13g2_o21ai_1
XFILLER_10_289 VPWR VGND sg13g2_fill_2
Xhold290 _0020_ VPWR VGND net837 sg13g2_dlygate4sd3_1
X_3225__218 VPWR VGND net218 sg13g2_tiehi
X_2521_ _0652_ net969 _1291_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_109 VPWR VGND sg13g2_fill_1
X_2452_ _0561_ _0581_ _0595_ VPWR VGND sg13g2_nor2_1
X_2383_ net545 VPWR _0527_ VGND _0494_ _0526_ sg13g2_o21ai_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_36_186 VPWR VGND sg13g2_fill_1
X_3004_ net116 VGND VPWR net776 controller.inst_mem.mem_data\[108\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_2719_ VPWR VGND _0821_ net447 net449 net707 _0822_ net480 sg13g2_a221oi_1
XFILLER_47_429 VPWR VGND sg13g2_decap_8
XFILLER_42_178 VPWR VGND sg13g2_fill_2
XFILLER_46_462 VPWR VGND sg13g2_decap_8
X_3208__71 VPWR VGND net71 sg13g2_tiehi
X_1952_ _1297_ _1298_ _1299_ VPWR VGND sg13g2_nor2b_1
X_1883_ _1224_ _1228_ _1219_ _1234_ VPWR VGND _1233_ sg13g2_nand4_1
XFILLER_44_0 VPWR VGND sg13g2_fill_1
X_2504_ VPWR VGND controller.alu_buffer.buffer\[10\] net463 net483 controller.alu_buffer.buffer\[8\]
+ _0638_ net472 sg13g2_a221oi_1
X_2435_ _0575_ _0576_ _0574_ _0578_ VPWR VGND _0577_ sg13g2_nand4_1
XFILLER_37_440 VPWR VGND sg13g2_decap_8
X_3144__81 VPWR VGND net81 sg13g2_tiehi
X_2366_ _0510_ VPWR _0511_ VGND net720 net491 sg13g2_o21ai_1
X_2297_ net531 _1206_ _1221_ _0443_ VPWR VGND sg13g2_nor3_1
XFILLER_20_373 VPWR VGND sg13g2_fill_2
XFILLER_46_42 VPWR VGND sg13g2_fill_1
XFILLER_43_443 VPWR VGND sg13g2_decap_8
XFILLER_15_112 VPWR VGND sg13g2_fill_2
X_2220_ VGND VPWR _1090_ net549 _0126_ _0385_ sg13g2_a21oi_1
X_2151_ net652 VPWR _0351_ VGND net810 net600 sg13g2_o21ai_1
X_2082_ VGND VPWR _1159_ net562 _0057_ _0316_ sg13g2_a21oi_1
X_2984_ net156 VGND VPWR _0007_ controller.inst_mem.mem_data\[88\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_1935_ net18 _1281_ _1282_ VPWR VGND sg13g2_nand2_1
X_1797_ VPWR _1148_ net735 VGND sg13g2_inv_1
X_1866_ controller.inst_mem.addr\[2\] _1216_ _1217_ VPWR VGND sg13g2_and2_1
X_2418_ VGND VPWR _0560_ _0561_ _0553_ _0546_ sg13g2_a21oi_2
XFILLER_29_226 VPWR VGND sg13g2_fill_1
X_2349_ _0495_ net524 controller.extended_jump_target\[0\] net499 controller.inst_mem.mem_data\[104\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_16_34 VPWR VGND sg13g2_fill_2
XFILLER_32_88 VPWR VGND sg13g2_fill_1
XFILLER_31_479 VPWR VGND sg13g2_fill_1
X_1651_ VPWR _1002_ net765 VGND sg13g2_inv_1
X_1720_ VPWR _1071_ net751 VGND sg13g2_inv_1
Xhold108 controller.inst_mem.mem_data\[136\] VPWR VGND net435 sg13g2_dlygate4sd3_1
XFILLER_7_196 VPWR VGND sg13g2_fill_1
Xhold119 controller.inst_mem.mem_data\[126\] VPWR VGND net666 sg13g2_dlygate4sd3_1
X_3252_ net67 VGND VPWR _0275_ controller.inst_mem.mem_data\[67\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3183_ net220 VGND VPWR net905 controller.counter2.counter_1\[14\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
X_2065_ net643 VPWR _0308_ VGND controller.inst_mem.mem_data\[130\] net585 sg13g2_o21ai_1
X_2203_ net649 VPWR _0377_ VGND controller.inst_mem.mem_data\[199\] net596 sg13g2_o21ai_1
X_2134_ VGND VPWR _1133_ net565 _0083_ _0342_ sg13g2_a21oi_1
X_2967_ net653 VPWR _0975_ VGND controller.inst_mem.mem_data\[76\] net601 sg13g2_o21ai_1
X_1849_ VPWR _1200_ net739 VGND sg13g2_inv_1
X_2898_ VGND VPWR _1020_ net554 _0249_ _0940_ sg13g2_a21oi_1
X_1918_ _1267_ _1261_ net917 _1256_ _1242_ VPWR VGND sg13g2_a22oi_1
XFILLER_45_505 VPWR VGND sg13g2_fill_2
X_3069__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_17_229 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_20_clk clknet_3_7__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_4_111 VPWR VGND sg13g2_fill_1
XFILLER_48_365 VPWR VGND sg13g2_decap_8
X_3200__135 VPWR VGND net135 sg13g2_tiehi
X_2821_ net636 VPWR _0902_ VGND controller.const_data\[3\] net570 sg13g2_o21ai_1
XFILLER_31_210 VPWR VGND sg13g2_fill_2
X_2683_ net448 VPWR _0794_ VGND _0409_ _0793_ sg13g2_o21ai_1
X_2752_ net452 _0847_ _0848_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_11_clk clknet_3_3__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_1703_ VPWR _1054_ net715 VGND sg13g2_inv_1
X_1634_ VPWR _0985_ net792 VGND sg13g2_inv_1
X_3235_ net107 VGND VPWR _0258_ controller.inst_mem.mem_data\[50\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_3166_ net288 VGND VPWR net900 controller.counter2.counter_0\[13\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
X_2048_ VGND VPWR _1176_ net618 _0040_ _0299_ sg13g2_a21oi_1
X_2117_ net630 VPWR _0334_ VGND controller.inst_mem.mem_data\[156\] net559 sg13g2_o21ai_1
X_3097_ net219 VGND VPWR net845 controller.extended_jump_target\[1\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
Xclkbuf_leaf_0_clk clknet_3_1__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
X_3020_ net84 VGND VPWR net743 controller.inst_mem.mem_data\[124\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_2804_ _0890_ _0884_ net904 VPWR VGND sg13g2_nand2b_1
X_2735_ net892 net915 _0834_ VPWR VGND sg13g2_xor2_1
X_2666_ VGND VPWR _0778_ _0779_ _0177_ _0780_ sg13g2_a21oi_1
X_2597_ VGND VPWR _1267_ _1268_ _0175_ _0503_ sg13g2_a21oi_1
XFILLER_39_184 VPWR VGND sg13g2_fill_2
X_3149_ net61 VGND VPWR net914 controller.alu_buffer.buffer\[23\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_3218_ net274 VGND VPWR _0241_ controller.inst_mem.mem_data\[33\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
Xhold291 controller.const_data\[3\] VPWR VGND net838 sg13g2_dlygate4sd3_1
XFILLER_2_412 VPWR VGND sg13g2_fill_2
Xhold280 _0286_ VPWR VGND net827 sg13g2_dlygate4sd3_1
X_2520_ controller.alu_buffer.buffer\[12\] _1291_ _0651_ VPWR VGND sg13g2_nor2_1
X_2451_ _0594_ _0590_ _0593_ VPWR VGND sg13g2_xnor2_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
X_3003_ net118 VGND VPWR net417 controller.inst_mem.mem_data\[107\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_2382_ _0525_ VPWR _0526_ VGND net486 _0523_ sg13g2_o21ai_1
X_2718_ _0821_ _0820_ _0417_ VPWR VGND sg13g2_nand2b_1
X_2649_ VGND VPWR _0485_ _0765_ _0764_ _0757_ sg13g2_a21oi_2
XFILLER_47_408 VPWR VGND sg13g2_decap_8
XFILLER_27_132 VPWR VGND sg13g2_fill_2
XFILLER_4_0 VPWR VGND sg13g2_fill_2
X_3051__311 VPWR VGND net311 sg13g2_tiehi
Xfanout590 net591 net590 VPWR VGND sg13g2_buf_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
X_1951_ controller.alu_buffer.buffer\[23\] controller.alu_buffer.buffer\[22\] controller.alu_buffer.buffer\[21\]
+ _1298_ VPWR VGND sg13g2_nor3_1
X_1882_ VPWR VGND controller.inst_mem.mem_data\[135\] net514 net519 controller.inst_mem.extended_word\[7\]
+ _1233_ net523 sg13g2_a221oi_1
XFILLER_37_0 VPWR VGND sg13g2_fill_2
X_2503_ VGND VPWR _0633_ _0636_ _0157_ _0637_ sg13g2_a21oi_1
X_2434_ _0577_ net496 controller.inst_mem.mem_data\[95\] net504 controller.inst_mem.mem_data\[191\]
+ VPWR VGND sg13g2_a22oi_1
X_2365_ _0507_ _0508_ _0506_ _0510_ VPWR VGND _0509_ sg13g2_nand4_1
X_2296_ net533 net536 net532 _0442_ VPWR VGND controller.extended_cond.opcode\[1\]
+ sg13g2_nand4_1
XFILLER_37_496 VPWR VGND sg13g2_decap_8
XFILLER_4_507 VPWR VGND sg13g2_fill_1
XFILLER_43_422 VPWR VGND sg13g2_decap_8
X_3261__238 VPWR VGND net238 sg13g2_tiehi
XFILLER_43_499 VPWR VGND sg13g2_decap_8
X_3079__255 VPWR VGND net255 sg13g2_tiehi
X_2081_ net632 VPWR _0316_ VGND controller.inst_mem.mem_data\[138\] net562 sg13g2_o21ai_1
X_2150_ VGND VPWR _1125_ net601 _0091_ _0350_ sg13g2_a21oi_1
X_3203__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_34_499 VPWR VGND sg13g2_decap_8
X_1934_ _1282_ _1279_ _1257_ _1258_ controller.alu_buffer.buffer\[3\] VPWR VGND sg13g2_a22oi_1
X_2983_ net158 VGND VPWR net785 controller.inst_mem.mem_data\[87\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_1796_ VPWR _1147_ net361 VGND sg13g2_inv_1
X_1865_ net534 net535 _1216_ VPWR VGND sg13g2_nor2b_1
X_2417_ _0559_ _0475_ _0485_ _0560_ VPWR VGND sg13g2_a21o_1
X_2348_ _0494_ _0486_ _0493_ VPWR VGND sg13g2_nand2_2
X_2279_ controller.extended_state\[0\] net535 _0425_ VPWR VGND sg13g2_xor2_1
XFILLER_40_469 VPWR VGND sg13g2_decap_8
XFILLER_32_78 VPWR VGND sg13g2_fill_1
X_1650_ VPWR _1001_ net809 VGND sg13g2_inv_1
Xhold109 controller.inst_mem.mem_data\[147\] VPWR VGND net436 sg13g2_dlygate4sd3_1
X_3182_ net224 VGND VPWR net927 controller.counter2.counter_1\[13\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
XFILLER_3_370 VPWR VGND sg13g2_fill_1
X_2202_ VGND VPWR _1099_ net599 _0117_ _0376_ sg13g2_a21oi_1
X_3251_ net99 VGND VPWR net375 controller.inst_mem.mem_data\[66\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_2064_ VGND VPWR _1168_ net586 _0048_ _0307_ sg13g2_a21oi_1
X_2133_ net633 VPWR _0342_ VGND net714 net565 sg13g2_o21ai_1
X_1917_ net16 _1265_ _1266_ VPWR VGND sg13g2_nand2_1
X_2897_ net635 VPWR _0940_ VGND controller.inst_mem.mem_data\[41\] net554 sg13g2_o21ai_1
X_2966_ VGND VPWR _0986_ net620 _0283_ _0974_ sg13g2_a21oi_1
X_1848_ VPWR _1199_ net421 VGND sg13g2_inv_1
X_1779_ VPWR _1130_ net425 VGND sg13g2_inv_1
XFILLER_25_252 VPWR VGND sg13g2_fill_2
X_2820_ VGND VPWR _1059_ net570 _0210_ _0901_ sg13g2_a21oi_1
X_2751_ _1270_ net903 _0847_ VPWR VGND sg13g2_xor2_1
X_2682_ _0408_ net938 _0793_ VPWR VGND sg13g2_nor2b_1
X_1702_ VPWR _1053_ net824 VGND sg13g2_inv_1
X_1633_ VPWR _0984_ net835 VGND sg13g2_inv_1
X_3165_ net292 VGND VPWR _0188_ controller.counter2.counter_0\[12\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
X_3234_ net123 VGND VPWR net408 controller.inst_mem.mem_data\[49\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_2047_ net662 VPWR _0299_ VGND net737 net621 sg13g2_o21ai_1
X_2116_ VGND VPWR _1142_ net581 _0074_ _0333_ sg13g2_a21oi_1
X_3096_ net221 VGND VPWR net830 controller.extended_jump_target\[0\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
X_2949_ net632 VPWR _0966_ VGND net767 net563 sg13g2_o21ai_1
XFILLER_1_137 VPWR VGND sg13g2_fill_1
Xhold440 _0148_ VPWR VGND net987 sg13g2_dlygate4sd3_1
XFILLER_38_33 VPWR VGND sg13g2_fill_2
X_3262__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_48_141 VPWR VGND sg13g2_fill_1
X_2734_ VGND VPWR net475 _0832_ _0192_ _0833_ sg13g2_a21oi_1
X_2803_ VGND VPWR net475 _0888_ _0205_ _0889_ sg13g2_a21oi_1
X_2665_ net540 VPWR _0780_ VGND net930 net444 sg13g2_o21ai_1
X_2596_ VGND VPWR _1265_ _1266_ _0174_ _0503_ sg13g2_a21oi_1
X_3148_ net65 VGND VPWR net957 controller.alu_buffer.buffer\[22\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_3217_ net282 VGND VPWR _0240_ controller.inst_mem.mem_data\[32\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_3079_ net255 VGND VPWR _0102_ controller.inst_mem.mem_data\[183\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
Xhold292 controller.inst_mem.mem_data\[119\] VPWR VGND net839 sg13g2_dlygate4sd3_1
Xhold270 _0019_ VPWR VGND net817 sg13g2_dlygate4sd3_1
Xhold281 controller.inst_mem.mem_data\[110\] VPWR VGND net828 sg13g2_dlygate4sd3_1
X_2450_ _0593_ _0591_ _0592_ VPWR VGND sg13g2_xnor2_1
X_2381_ _0525_ _0517_ _0524_ VPWR VGND sg13g2_nand2b_1
XFILLER_49_494 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[5] net5 VPWR VGND sg13g2_buf_1
X_3089__235 VPWR VGND net235 sg13g2_tiehi
X_3002_ net120 VGND VPWR _0025_ controller.inst_mem.mem_data\[106\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
X_2717_ net899 VPWR _0820_ VGND controller.counter2.counter_0\[12\] _0415_ sg13g2_o21ai_1
X_2648_ _0758_ _0763_ _0475_ _0764_ VPWR VGND sg13g2_nand3_1
X_2579_ _0695_ net956 _0700_ VPWR VGND sg13g2_xor2_1
X_3217__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_46_420 VPWR VGND sg13g2_decap_8
Xfanout580 net624 net580 VPWR VGND sg13g2_buf_8
Xfanout591 net605 net591 VPWR VGND sg13g2_buf_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
X_3229__186 VPWR VGND net186 sg13g2_tiehi
X_1950_ _1297_ _1296_ controller.alu_buffer.buffer\[20\] VPWR VGND sg13g2_nand2b_1
X_2502_ net539 VPWR _0637_ VGND net973 net460 sg13g2_o21ai_1
X_1881_ _1232_ _1068_ net520 VPWR VGND sg13g2_nand2_1
X_2433_ _0576_ net525 controller.extended_then_action\[3\] net500 controller.inst_mem.mem_data\[119\]
+ VPWR VGND sg13g2_a22oi_1
X_2364_ _0509_ _0479_ controller.inst_mem.mem_data\[129\] net524 controller.extended_jump_target\[1\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_49_280 VPWR VGND sg13g2_fill_1
XFILLER_37_475 VPWR VGND sg13g2_decap_8
X_2295_ _1110_ _1223_ _0441_ VPWR VGND sg13g2_nor2_1
XANTENNA_10 VPWR VGND uio_in[5] sg13g2_antennanp
XFILLER_21_58 VPWR VGND sg13g2_fill_2
XFILLER_43_478 VPWR VGND sg13g2_decap_8
X_2080_ VGND VPWR _1160_ net558 _0056_ _0315_ sg13g2_a21oi_1
XFILLER_34_478 VPWR VGND sg13g2_decap_8
X_2982_ net160 VGND VPWR _0005_ controller.inst_mem.mem_data\[86\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_1933_ _1281_ controller.alu_buffer.buffer\[19\] _1260_ VPWR VGND sg13g2_nand2_1
X_3039__46 VPWR VGND net46 sg13g2_tiehi
X_1864_ VPWR _1215_ net705 VGND sg13g2_inv_1
X_1795_ VPWR _1146_ net357 VGND sg13g2_inv_1
X_2416_ _0558_ VPWR _0559_ VGND controller.inst_mem.mem_data\[49\] net491 sg13g2_o21ai_1
X_2347_ net486 _0491_ net488 _0493_ VPWR VGND _0492_ sg13g2_nand4_1
X_2278_ controller.extended_state\[1\] net534 _0424_ VPWR VGND sg13g2_xor2_1
XFILLER_40_448 VPWR VGND sg13g2_decap_8
XFILLER_32_35 VPWR VGND sg13g2_fill_2
XFILLER_4_316 VPWR VGND sg13g2_fill_1
X_3115__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_43_286 VPWR VGND sg13g2_fill_2
X_3181_ net228 VGND VPWR _0204_ controller.counter2.counter_1\[12\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_2201_ net652 VPWR _0376_ VGND controller.inst_mem.mem_data\[198\] net599 sg13g2_o21ai_1
X_3250_ net131 VGND VPWR net329 controller.inst_mem.mem_data\[65\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_2132_ VGND VPWR _1134_ net563 _0082_ _0341_ sg13g2_a21oi_1
X_2063_ net643 VPWR _0307_ VGND net340 net587 sg13g2_o21ai_1
XFILLER_19_250 VPWR VGND sg13g2_fill_2
X_1847_ VPWR _1198_ net708 VGND sg13g2_inv_1
X_2896_ VGND VPWR _1021_ net547 _0248_ _0939_ sg13g2_a21oi_1
X_2965_ net651 VPWR _0974_ VGND controller.inst_mem.mem_data\[75\] net601 sg13g2_o21ai_1
X_1916_ _1266_ _1260_ controller.alu_buffer.buffer\[17\] _1258_ net530 VPWR VGND sg13g2_a22oi_1
X_1778_ VPWR _1129_ net350 VGND sg13g2_inv_1
XFILLER_45_507 VPWR VGND sg13g2_fill_1
XFILLER_36_507 VPWR VGND sg13g2_fill_1
X_3048__317 VPWR VGND net317 sg13g2_tiehi
XFILLER_16_231 VPWR VGND sg13g2_fill_1
X_2681_ VGND VPWR _0790_ _0791_ _0180_ _0792_ sg13g2_a21oi_1
X_1701_ VPWR _1052_ net788 VGND sg13g2_inv_1
X_2750_ VGND VPWR net477 _0845_ _0195_ _0846_ sg13g2_a21oi_1
X_1632_ VPWR _0983_ net826 VGND sg13g2_inv_1
X_3164_ net296 VGND VPWR net898 controller.counter2.counter_0\[11\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
X_3233_ net139 VGND VPWR _0256_ controller.inst_mem.mem_data\[48\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_2115_ net642 VPWR _0333_ VGND net703 net581 sg13g2_o21ai_1
X_3095_ net223 VGND VPWR net756 controller.inst_mem.mem_data\[199\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_2046_ VGND VPWR _1177_ net617 _0039_ _0298_ sg13g2_a21oi_1
X_3099__215 VPWR VGND net215 sg13g2_tiehi
X_2948_ VGND VPWR _0995_ net562 _0274_ _0965_ sg13g2_a21oi_1
X_2879_ net646 VPWR _0931_ VGND net777 net590 sg13g2_o21ai_1
Xhold430 controller.alu_buffer.buffer\[3\] VPWR VGND net977 sg13g2_dlygate4sd3_1
XFILLER_18_507 VPWR VGND sg13g2_fill_1
X_3014__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_5_444 VPWR VGND sg13g2_fill_1
XFILLER_44_381 VPWR VGND sg13g2_fill_1
X_2664_ VPWR VGND net8 net446 _0774_ net695 _0779_ net479 sg13g2_a221oi_1
X_2733_ net544 VPWR _0833_ VGND net892 net475 sg13g2_o21ai_1
X_2802_ net544 VPWR _0889_ VGND net926 net474 sg13g2_o21ai_1
X_2595_ net15 net537 _0173_ VPWR VGND sg13g2_and2_1
X_3216_ net290 VGND VPWR net690 controller.const_data\[31\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_27_304 VPWR VGND sg13g2_fill_1
X_3147_ net69 VGND VPWR _0170_ controller.alu_buffer.buffer\[21\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
X_3078_ net257 VGND VPWR net849 controller.inst_mem.mem_data\[182\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_2029_ net628 VPWR _0290_ VGND controller.inst_mem.mem_data\[112\] net552 sg13g2_o21ai_1
Xhold271 controller.const_data\[26\] VPWR VGND net818 sg13g2_dlygate4sd3_1
Xhold260 controller.inst_mem.mem_data\[60\] VPWR VGND net807 sg13g2_dlygate4sd3_1
Xhold293 controller.const_data\[22\] VPWR VGND net840 sg13g2_dlygate4sd3_1
Xhold282 controller.inst_mem.mem_data\[199\] VPWR VGND net829 sg13g2_dlygate4sd3_1
XFILLER_18_304 VPWR VGND sg13g2_fill_1
X_2380_ net486 VPWR _0524_ VGND controller.extended_jump_target\[2\] net488 sg13g2_o21ai_1
XFILLER_49_473 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[6] net6 VPWR VGND sg13g2_buf_1
X_3001_ net122 VGND VPWR net389 controller.inst_mem.mem_data\[105\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
XFILLER_32_384 VPWR VGND sg13g2_fill_1
X_2716_ VGND VPWR net445 _0818_ _0188_ _0819_ sg13g2_a21oi_1
X_2647_ _0761_ _0762_ _0760_ _0763_ VPWR VGND sg13g2_nand3_1
X_2578_ _0699_ _0695_ controller.alu_buffer.buffer\[22\] VPWR VGND sg13g2_nand2b_1
XFILLER_27_189 VPWR VGND sg13g2_fill_2
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
X_3153__51 VPWR VGND net51 sg13g2_tiehi
Xfanout570 net571 net570 VPWR VGND sg13g2_buf_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
Xfanout581 net584 net581 VPWR VGND sg13g2_buf_8
Xfanout592 net594 net592 VPWR VGND sg13g2_buf_8
XFILLER_18_189 VPWR VGND sg13g2_fill_2
X_1880_ net532 net533 net536 _1231_ VPWR VGND sg13g2_nor3_2
X_2501_ _0636_ _0635_ net468 net457 net14 VPWR VGND sg13g2_a22oi_1
X_2363_ _0508_ net499 controller.inst_mem.mem_data\[105\] net503 controller.inst_mem.mem_data\[177\]
+ VPWR VGND sg13g2_a22oi_1
X_2294_ net844 net488 _0440_ VPWR VGND sg13g2_nor2_1
X_2432_ VPWR VGND controller.inst_mem.mem_data\[143\] net518 net520 controller.inst_mem.mem_data\[167\]
+ _0575_ net512 sg13g2_a221oi_1
XFILLER_37_454 VPWR VGND sg13g2_decap_8
XANTENNA_11 VPWR VGND uio_in[6] sg13g2_antennanp
XFILLER_20_332 VPWR VGND sg13g2_fill_2
XFILLER_43_457 VPWR VGND sg13g2_decap_8
XFILLER_11_376 VPWR VGND sg13g2_fill_2
XFILLER_34_457 VPWR VGND sg13g2_decap_8
X_1932_ _1276_ _1278_ _1274_ _1280_ VPWR VGND sg13g2_nand3_1
X_2981_ net162 VGND VPWR net725 controller.inst_mem.mem_data\[85\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_1863_ VPWR _1214_ net677 VGND sg13g2_inv_1
X_2415_ _0555_ _0556_ _0554_ _0558_ VPWR VGND _0557_ sg13g2_nand4_1
X_1794_ VPWR _1145_ net797 VGND sg13g2_inv_1
XFILLER_37_240 VPWR VGND sg13g2_fill_1
X_2346_ _0492_ _1025_ net517 VPWR VGND sg13g2_nand2_1
X_2277_ controller.extended_state\[2\] net532 _0423_ VPWR VGND sg13g2_xor2_1
XFILLER_40_416 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_32_clk clknet_3_4__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_48_505 VPWR VGND sg13g2_fill_2
XFILLER_0_501 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_3_4__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
X_3233__139 VPWR VGND net139 sg13g2_tiehi
X_3180_ net232 VGND VPWR net884 controller.counter2.counter_1\[11\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_2062_ VGND VPWR _1169_ net592 _0047_ _0306_ sg13g2_a21oi_1
X_2200_ VGND VPWR _1100_ net599 _0116_ _0375_ sg13g2_a21oi_1
X_2131_ net632 VPWR _0341_ VGND net732 net563 sg13g2_o21ai_1
XFILLER_34_265 VPWR VGND sg13g2_fill_2
XFILLER_34_232 VPWR VGND sg13g2_fill_1
X_2964_ VGND VPWR _0987_ net619 _0282_ _0973_ sg13g2_a21oi_1
X_3244__246 VPWR VGND net246 sg13g2_tiehi
XFILLER_22_416 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_14_clk clknet_3_6__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
XFILLER_30_471 VPWR VGND sg13g2_fill_1
X_1846_ VPWR _1197_ net816 VGND sg13g2_inv_1
X_2895_ net627 VPWR _0939_ VGND net722 net547 sg13g2_o21ai_1
X_1777_ VPWR _1128_ net336 VGND sg13g2_inv_1
X_1915_ _1265_ _1261_ net940 _1256_ _1236_ VPWR VGND sg13g2_a22oi_1
X_2329_ VGND VPWR _0475_ _0473_ _0469_ sg13g2_or2_1
X_3026__72 VPWR VGND net72 sg13g2_tiehi
XFILLER_13_405 VPWR VGND sg13g2_fill_2
X_3041__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_48_379 VPWR VGND sg13g2_decap_8
X_2680_ net540 VPWR _0792_ VGND net944 net444 sg13g2_o21ai_1
X_1700_ VPWR _1051_ net390 VGND sg13g2_inv_1
X_1631_ VPWR _0982_ net874 VGND sg13g2_inv_1
X_3239__326 VPWR VGND net326 sg13g2_tiehi
X_3232_ net155 VGND VPWR _0255_ controller.inst_mem.mem_data\[47\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_3_clk clknet_3_2__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ net300 VGND VPWR net925 controller.counter2.counter_0\[10\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
X_2045_ net662 VPWR _0298_ VGND net760 net617 sg13g2_o21ai_1
X_2114_ VGND VPWR _1143_ net585 _0073_ _0332_ sg13g2_a21oi_1
X_3094_ net225 VGND VPWR net712 controller.inst_mem.mem_data\[198\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_2947_ net632 VPWR _0965_ VGND controller.inst_mem.mem_data\[66\] net562 sg13g2_o21ai_1
Xhold420 controller.alu_buffer.buffer\[8\] VPWR VGND net967 sg13g2_dlygate4sd3_1
X_2878_ VGND VPWR _1030_ net574 _0239_ _0930_ sg13g2_a21oi_1
Xhold431 controller.inst_mem.addr\[1\] VPWR VGND net978 sg13g2_dlygate4sd3_1
X_1829_ VPWR _1180_ net673 VGND sg13g2_inv_1
X_2801_ VGND VPWR net440 net450 _0888_ _0887_ sg13g2_a21oi_1
X_2732_ VGND VPWR net418 net451 _0832_ _0831_ sg13g2_a21oi_1
X_2663_ net448 VPWR _0778_ VGND _0405_ _0777_ sg13g2_o21ai_1
X_2594_ VGND VPWR net459 _0712_ _0172_ _0713_ sg13g2_a21oi_1
X_3215_ net298 VGND VPWR net441 controller.const_data\[30\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_39_110 VPWR VGND sg13g2_fill_1
X_3077_ net259 VGND VPWR net399 controller.inst_mem.mem_data\[181\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_2028_ VGND VPWR _1186_ net548 _0030_ _0289_ sg13g2_a21oi_1
X_3146_ net73 VGND VPWR net949 controller.alu_buffer.buffer\[20\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
Xhold261 _0269_ VPWR VGND net808 sg13g2_dlygate4sd3_1
Xhold294 controller.inst_mem.mem_data\[153\] VPWR VGND net841 sg13g2_dlygate4sd3_1
Xhold283 _0119_ VPWR VGND net830 sg13g2_dlygate4sd3_1
Xhold250 controller.inst_mem.mem_data\[151\] VPWR VGND net797 sg13g2_dlygate4sd3_1
Xhold272 controller.inst_mem.mem_data\[115\] VPWR VGND net819 sg13g2_dlygate4sd3_1
XFILLER_45_146 VPWR VGND sg13g2_fill_2
XFILLER_49_452 VPWR VGND sg13g2_decap_8
Xinput7 uio_in[0] net7 VPWR VGND sg13g2_buf_1
X_3000_ net124 VGND VPWR _0023_ controller.inst_mem.mem_data\[104\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
X_2715_ net541 VPWR _0819_ VGND net916 net445 sg13g2_o21ai_1
X_2577_ VGND VPWR _0694_ _0697_ _0170_ _0698_ sg13g2_a21oi_1
X_2646_ VPWR VGND controller.inst_mem.mem_data\[116\] _0759_ net501 controller.inst_mem.mem_data\[164\]
+ _0762_ net513 sg13g2_a221oi_1
X_3129_ net141 VGND VPWR _0152_ controller.alu_buffer.buffer\[2\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_7_507 VPWR VGND sg13g2_fill_1
Xfanout560 net561 net560 VPWR VGND sg13g2_buf_1
XFILLER_46_455 VPWR VGND sg13g2_decap_8
Xfanout571 net580 net571 VPWR VGND sg13g2_buf_8
Xfanout582 net584 net582 VPWR VGND sg13g2_buf_8
Xfanout593 net594 net593 VPWR VGND sg13g2_buf_8
X_2500_ _0635_ _1287_ _0634_ VPWR VGND sg13g2_nand2_1
X_2431_ _0574_ controller.inst_mem.mem_data\[71\] net508 VPWR VGND sg13g2_nand2_1
X_2293_ VGND VPWR _0439_ net489 _0422_ sg13g2_or2_1
XFILLER_2_84 VPWR VGND sg13g2_fill_1
X_2362_ _0507_ net495 controller.inst_mem.mem_data\[81\] net511 controller.inst_mem.mem_data\[153\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_24_149 VPWR VGND sg13g2_fill_2
XANTENNA_12 VPWR VGND uio_in[7] sg13g2_antennanp
XFILLER_20_366 VPWR VGND sg13g2_fill_2
X_2629_ _0744_ VPWR _0745_ VGND controller.inst_mem.mem_data\[46\] net492 sg13g2_o21ai_1
XFILLER_28_444 VPWR VGND sg13g2_fill_1
XFILLER_43_436 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_fill_2
X_2980_ net164 VGND VPWR _0003_ controller.inst_mem.mem_data\[84\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
Xinput10 uio_in[3] net10 VPWR VGND sg13g2_buf_1
XFILLER_42_491 VPWR VGND sg13g2_decap_8
X_1931_ _1277_ _1278_ _1279_ VPWR VGND sg13g2_nor2b_2
X_1793_ VPWR _1144_ net771 VGND sg13g2_inv_1
X_1862_ VPWR _1213_ net778 VGND sg13g2_inv_1
X_2414_ VPWR VGND controller.inst_mem.mem_data\[145\] net518 net520 controller.inst_mem.mem_data\[97\]
+ _0557_ net495 sg13g2_a221oi_1
XFILLER_6_370 VPWR VGND sg13g2_fill_2
X_2276_ _0419_ _0421_ _0422_ VPWR VGND sg13g2_and2_1
X_2345_ _0488_ _0489_ _0487_ _0491_ VPWR VGND _0490_ sg13g2_nand4_1
X_2061_ net648 VPWR _0306_ VGND net773 net592 sg13g2_o21ai_1
X_2130_ VGND VPWR _1135_ net554 _0081_ _0340_ sg13g2_a21oi_1
X_2963_ net661 VPWR _0973_ VGND controller.inst_mem.mem_data\[74\] net619 sg13g2_o21ai_1
XFILLER_15_480 VPWR VGND sg13g2_fill_1
X_1914_ _1264_ VPWR net15 VGND _1067_ _1259_ sg13g2_o21ai_1
XFILLER_22_439 VPWR VGND sg13g2_fill_2
X_1845_ VPWR _1196_ net836 VGND sg13g2_inv_1
X_2894_ VGND VPWR _1022_ net551 _0247_ _0938_ sg13g2_a21oi_1
X_1776_ VPWR _1127_ net753 VGND sg13g2_inv_1
X_2328_ _0469_ _0473_ _0474_ VPWR VGND sg13g2_nor2_1
X_2259_ net930 controller.counter2.counter_0\[0\] _0405_ VPWR VGND sg13g2_nor2_1
XFILLER_27_59 VPWR VGND sg13g2_fill_2
X_2980__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_0_310 VPWR VGND sg13g2_fill_1
X_1630_ VPWR _0981_ net691 VGND sg13g2_inv_1
X_3162_ net304 VGND VPWR net887 controller.counter2.counter_0\[9\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
X_3231_ net170 VGND VPWR net665 controller.inst_mem.mem_data\[46\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
XFILLER_47_380 VPWR VGND sg13g2_decap_8
X_2044_ VGND VPWR _1178_ net609 _0038_ _0297_ sg13g2_a21oi_1
X_2113_ net643 VPWR _0332_ VGND net823 net585 sg13g2_o21ai_1
X_3093_ net227 VGND VPWR _0116_ controller.inst_mem.mem_data\[197\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_2877_ net638 VPWR _0930_ VGND controller.const_data\[31\] net574 sg13g2_o21ai_1
X_2946_ VGND VPWR _0996_ net552 _0273_ _0964_ sg13g2_a21oi_1
Xhold421 _0149_ VPWR VGND net968 sg13g2_dlygate4sd3_1
Xhold410 _0171_ VPWR VGND net957 sg13g2_dlygate4sd3_1
Xhold432 _0147_ VPWR VGND net979 sg13g2_dlygate4sd3_1
X_1759_ VPWR _1110_ net814 VGND sg13g2_inv_1
X_1828_ VPWR _1179_ net779 VGND sg13g2_inv_1
XFILLER_13_258 VPWR VGND sg13g2_fill_1
X_2731_ net892 net451 _0831_ VPWR VGND sg13g2_nor2_1
X_2800_ net450 _0886_ _0887_ VPWR VGND sg13g2_nor2_1
X_2662_ net930 controller.counter2.counter_0\[0\] _0777_ VPWR VGND sg13g2_and2_1
X_2593_ net537 VPWR _0713_ VGND net913 net459 sg13g2_o21ai_1
X_3214_ net306 VGND VPWR _0237_ controller.const_data\[29\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3145_ net77 VGND VPWR net946 controller.alu_buffer.buffer\[19\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
X_2027_ net625 VPWR _0289_ VGND net730 net549 sg13g2_o21ai_1
X_3076_ net261 VGND VPWR _0099_ controller.inst_mem.mem_data\[180\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_2929_ net644 VPWR _0956_ VGND net426 net587 sg13g2_o21ai_1
Xhold273 controller.const_data\[23\] VPWR VGND net820 sg13g2_dlygate4sd3_1
Xhold284 controller.inst_mem.mem_data\[131\] VPWR VGND net831 sg13g2_dlygate4sd3_1
Xhold262 controller.inst_mem.mem_data\[59\] VPWR VGND net809 sg13g2_dlygate4sd3_1
Xhold295 controller.extended_jump_target\[2\] VPWR VGND net842 sg13g2_dlygate4sd3_1
Xhold251 controller.inst_mem.mem_data\[127\] VPWR VGND net798 sg13g2_dlygate4sd3_1
Xhold240 _0261_ VPWR VGND net787 sg13g2_dlygate4sd3_1
X_3264__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_41_320 VPWR VGND sg13g2_fill_1
XFILLER_26_372 VPWR VGND sg13g2_fill_1
XFILLER_49_431 VPWR VGND sg13g2_decap_8
Xinput8 uio_in[1] net8 VPWR VGND sg13g2_buf_1
X_2714_ _0818_ net449 _0817_ _0767_ net372 VPWR VGND sg13g2_a22oi_1
X_2645_ _0761_ net494 controller.inst_mem.mem_data\[92\] net509 controller.inst_mem.mem_data\[68\]
+ VPWR VGND sg13g2_a22oi_1
X_2576_ net537 VPWR _0698_ VGND net960 net458 sg13g2_o21ai_1
X_3128_ net145 VGND VPWR _0151_ controller.alu_buffer.buffer\[1\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_3059_ net295 VGND VPWR _0082_ controller.inst_mem.mem_data\[163\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
Xfanout572 net574 net572 VPWR VGND sg13g2_buf_8
Xfanout550 net553 net550 VPWR VGND sg13g2_buf_8
Xfanout583 net584 net583 VPWR VGND sg13g2_buf_1
Xfanout561 net568 net561 VPWR VGND sg13g2_buf_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
Xfanout594 net605 net594 VPWR VGND sg13g2_buf_8
XFILLER_25_92 VPWR VGND sg13g2_fill_1
XFILLER_14_342 VPWR VGND sg13g2_fill_1
X_2430_ _0564_ _0572_ net487 _0573_ VPWR VGND sg13g2_nand3_1
X_2361_ VGND VPWR controller.inst_mem.mem_data\[57\] net507 _0506_ net517 sg13g2_a21oi_1
X_2292_ _0426_ VPWR _0438_ VGND _0421_ _0437_ sg13g2_o21ai_1
XANTENNA_13 VPWR VGND ui_in[1] sg13g2_antennanp
XFILLER_37_489 VPWR VGND sg13g2_decap_8
X_3104__205 VPWR VGND net205 sg13g2_tiehi
X_2628_ _0742_ _0743_ _0740_ _0744_ VPWR VGND sg13g2_nand3_1
X_2559_ net537 VPWR _0684_ VGND net952 net458 sg13g2_o21ai_1
XFILLER_46_58 VPWR VGND sg13g2_fill_2
XFILLER_43_415 VPWR VGND sg13g2_decap_8
XFILLER_28_412 VPWR VGND sg13g2_fill_1
X_3005__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_23_183 VPWR VGND sg13g2_fill_2
X_2990__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_42_470 VPWR VGND sg13g2_decap_8
X_1930_ controller.counter2.counter_1\[15\] controller.counter2.counter_1\[14\] controller.counter2.counter_1\[13\]
+ controller.counter2.counter_1\[12\] _1278_ VPWR VGND sg13g2_nor4_1
Xinput11 uio_in[4] net11 VPWR VGND sg13g2_buf_1
X_1861_ VPWR _1212_ net724 VGND sg13g2_inv_1
X_1792_ VPWR _1143_ net841 VGND sg13g2_inv_1
X_2413_ _0556_ net525 controller.extended_then_action\[5\] net507 controller.inst_mem.mem_data\[73\]
+ VPWR VGND sg13g2_a22oi_1
X_2344_ VPWR VGND controller.inst_mem.mem_data\[131\] net517 net520 controller.inst_mem.mem_data\[107\]
+ _0490_ net498 sg13g2_a221oi_1
X_2275_ controller.extended_cond.opcode\[2\] controller.extended_cond.opcode\[1\]
+ controller.extended_cond.opcode\[0\] _0421_ VPWR VGND sg13g2_nor3_1
XFILLER_48_507 VPWR VGND sg13g2_fill_1
XFILLER_43_223 VPWR VGND sg13g2_fill_2
XFILLER_28_264 VPWR VGND sg13g2_fill_2
X_2060_ VGND VPWR _1170_ net596 _0046_ _0305_ sg13g2_a21oi_1
XFILLER_19_286 VPWR VGND sg13g2_fill_1
X_2962_ VGND VPWR _0988_ net616 _0281_ _0972_ sg13g2_a21oi_1
X_2893_ net626 VPWR _0938_ VGND net799 net547 sg13g2_o21ai_1
X_1913_ VGND VPWR net965 _1260_ _1264_ _1263_ sg13g2_a21oi_1
X_1844_ VPWR _1195_ net860 VGND sg13g2_inv_1
X_1775_ VPWR _1126_ net780 VGND sg13g2_inv_1
X_2327_ VPWR VGND _0472_ _0466_ _0471_ _0457_ _0473_ _0470_ sg13g2_a221oi_1
X_2258_ VGND VPWR _1071_ net588 _0145_ _0404_ sg13g2_a21oi_1
X_2189_ net662 VPWR _0370_ VGND controller.inst_mem.mem_data\[192\] net617 sg13g2_o21ai_1
XFILLER_25_267 VPWR VGND sg13g2_fill_1
X_3191__188 VPWR VGND net188 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_30 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_48_337 VPWR VGND sg13g2_fill_1
XFILLER_8_411 VPWR VGND sg13g2_fill_1
XFILLER_8_466 VPWR VGND sg13g2_fill_2
X_3161_ net308 VGND VPWR _0184_ controller.counter2.counter_0\[8\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_3230_ net178 VGND VPWR _0253_ controller.inst_mem.mem_data\[45\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_2112_ VGND VPWR _1144_ net586 _0072_ _0331_ sg13g2_a21oi_1
X_2043_ net656 VPWR _0297_ VGND controller.inst_mem.mem_data\[119\] net609 sg13g2_o21ai_1
X_3092_ net229 VGND VPWR net791 controller.inst_mem.mem_data\[196\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_2876_ VGND VPWR _1031_ net576 _0238_ _0929_ sg13g2_a21oi_1
X_1827_ VPWR _1178_ net768 VGND sg13g2_inv_1
X_2945_ net629 VPWR _0964_ VGND controller.inst_mem.mem_data\[65\] net552 sg13g2_o21ai_1
X_1689_ VPWR _1040_ net736 VGND sg13g2_inv_1
Xhold400 controller.counter2.counter_0\[0\] VPWR VGND net947 sg13g2_dlygate4sd3_1
Xhold433 controller.alu_buffer.buffer\[5\] VPWR VGND net980 sg13g2_dlygate4sd3_1
Xhold422 controller.alu_buffer.buffer\[12\] VPWR VGND net969 sg13g2_dlygate4sd3_1
Xhold411 controller.alu_buffer.buffer\[17\] VPWR VGND net958 sg13g2_dlygate4sd3_1
X_1758_ VPWR _1109_ net834 VGND sg13g2_inv_1
X_3112__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_41_502 VPWR VGND sg13g2_decap_4
XFILLER_32_502 VPWR VGND sg13g2_decap_4
X_2661_ VGND VPWR _0771_ _0775_ _0176_ _0776_ sg13g2_a21oi_1
X_2730_ VGND VPWR _0830_ _0765_ net480 sg13g2_or2_1
X_2592_ _0711_ VPWR _0712_ VGND _0707_ _0710_ sg13g2_o21ai_1
X_3213_ net314 VGND VPWR net397 controller.const_data\[28\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3075_ net263 VGND VPWR _0098_ controller.inst_mem.mem_data\[179\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
X_3144_ net81 VGND VPWR net953 controller.alu_buffer.buffer\[18\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
X_2026_ VGND VPWR _1187_ net550 _0029_ _1339_ sg13g2_a21oi_1
X_2859_ net658 VPWR _0921_ VGND controller.const_data\[22\] net613 sg13g2_o21ai_1
X_2928_ VGND VPWR _1005_ net593 _0264_ _0955_ sg13g2_a21oi_1
Xhold241 controller.const_data\[8\] VPWR VGND net788 sg13g2_dlygate4sd3_1
Xhold285 controller.const_data\[2\] VPWR VGND net832 sg13g2_dlygate4sd3_1
Xhold274 controller.inst_mem.mem_data\[95\] VPWR VGND net821 sg13g2_dlygate4sd3_1
Xhold263 controller.inst_mem.mem_data\[173\] VPWR VGND net810 sg13g2_dlygate4sd3_1
Xhold230 controller.inst_mem.mem_data\[32\] VPWR VGND net777 sg13g2_dlygate4sd3_1
Xhold252 controller.inst_mem.mem_data\[39\] VPWR VGND net799 sg13g2_dlygate4sd3_1
Xhold296 controller.inst_mem.mem_data\[196\] VPWR VGND net843 sg13g2_dlygate4sd3_1
XFILLER_18_318 VPWR VGND sg13g2_fill_1
XFILLER_30_82 VPWR VGND sg13g2_fill_1
XFILLER_5_244 VPWR VGND sg13g2_fill_1
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
Xinput9 uio_in[2] net9 VPWR VGND sg13g2_buf_1
XFILLER_32_365 VPWR VGND sg13g2_fill_1
X_3065__283 VPWR VGND net283 sg13g2_tiehi
X_2713_ _0817_ net916 _0415_ VPWR VGND sg13g2_xnor2_1
X_2644_ _0760_ net526 controller.extended_then_action\[0\] net505 controller.inst_mem.mem_data\[188\]
+ VPWR VGND sg13g2_a22oi_1
X_2575_ _0697_ _0696_ net466 net455 net954 VPWR VGND sg13g2_a22oi_1
X_3127_ net149 VGND VPWR net972 controller.alu_buffer.buffer\[0\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_2
X_3058_ net297 VGND VPWR net339 controller.inst_mem.mem_data\[162\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_2009_ net649 VPWR _1331_ VGND controller.inst_mem.mem_data\[102\] net595 sg13g2_o21ai_1
X_2977__115 VPWR VGND net115 sg13g2_tiehi
Xfanout540 net541 net540 VPWR VGND sg13g2_buf_1
XFILLER_46_413 VPWR VGND sg13g2_decap_8
Xfanout573 net574 net573 VPWR VGND sg13g2_buf_1
Xfanout584 net591 net584 VPWR VGND sg13g2_buf_8
Xfanout595 net596 net595 VPWR VGND sg13g2_buf_8
Xfanout551 net553 net551 VPWR VGND sg13g2_buf_8
Xfanout562 net564 net562 VPWR VGND sg13g2_buf_8
X_2291_ VPWR VGND _1300_ _0435_ _0436_ _1280_ _0437_ _0420_ sg13g2_a221oi_1
X_2360_ _0505_ net534 net536 VPWR VGND sg13g2_xnor2_1
XFILLER_37_468 VPWR VGND sg13g2_decap_8
XANTENNA_14 VPWR VGND uio_in[3] sg13g2_antennanp
X_2627_ VPWR VGND controller.extended_then_action\[2\] _0741_ net525 controller.inst_mem.mem_data\[190\]
+ _0743_ net504 sg13g2_a221oi_1
X_2489_ _1285_ VPWR _0626_ VGND _1066_ _0622_ sg13g2_o21ai_1
X_2558_ _0683_ net455 controller.alu_buffer.buffer\[10\] net470 controller.alu_buffer.buffer\[17\]
+ VPWR VGND sg13g2_a22oi_1
X_3150__57 VPWR VGND net57 sg13g2_tiehi
Xclkbuf_leaf_35_clk clknet_3_1__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_11_40 VPWR VGND sg13g2_fill_2
XFILLER_46_210 VPWR VGND sg13g2_fill_2
XFILLER_19_424 VPWR VGND sg13g2_fill_2
X_3166__288 VPWR VGND net288 sg13g2_tiehi
X_1860_ VPWR _1211_ net796 VGND sg13g2_inv_1
Xclkbuf_leaf_26_clk clknet_3_5__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
Xinput12 uio_in[5] net12 VPWR VGND sg13g2_buf_1
X_1791_ VPWR _1142_ net823 VGND sg13g2_inv_1
X_2274_ controller.extended_cond.opcode\[2\] controller.extended_cond.opcode\[1\]
+ _0420_ VPWR VGND sg13g2_nor2_1
X_2412_ _0555_ net503 controller.inst_mem.mem_data\[193\] net511 controller.inst_mem.mem_data\[169\]
+ VPWR VGND sg13g2_a22oi_1
X_2343_ _0489_ net494 controller.inst_mem.mem_data\[83\] net510 controller.inst_mem.mem_data\[155\]
+ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_17_clk clknet_3_7__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_33_493 VPWR VGND sg13g2_decap_8
X_1989_ net633 VPWR _1321_ VGND controller.inst_mem.mem_data\[92\] net567 sg13g2_o21ai_1
X_3122__169 VPWR VGND net169 sg13g2_tiehi
X_2961_ net660 VPWR _0972_ VGND net346 net616 sg13g2_o21ai_1
X_1843_ VPWR _1194_ net865 VGND sg13g2_inv_1
X_2892_ VGND VPWR _1023_ net558 _0246_ _0937_ sg13g2_a21oi_1
X_1912_ _1255_ _1262_ _1263_ VPWR VGND sg13g2_nor2_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_1774_ VPWR _1125_ net744 VGND sg13g2_inv_1
Xclkbuf_leaf_6_clk clknet_3_2__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_6_191 VPWR VGND sg13g2_fill_2
X_2326_ VGND VPWR net4 _0448_ _0472_ _0457_ sg13g2_a21oi_1
X_2257_ net647 VPWR _0404_ VGND controller.extended_state\[2\] net588 sg13g2_o21ai_1
XFILLER_40_249 VPWR VGND sg13g2_fill_2
X_3259__83 VPWR VGND net83 sg13g2_tiehi
X_2188_ VGND VPWR _1106_ net609 _0110_ _0369_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_31 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_0_345 VPWR VGND sg13g2_fill_2
X_3160_ net312 VGND VPWR net880 controller.counter2.counter_0\[7\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
X_2042_ VGND VPWR _1179_ net606 _0037_ _0296_ sg13g2_a21oi_1
X_3091_ net231 VGND VPWR net401 controller.inst_mem.mem_data\[195\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_2
X_2111_ net643 VPWR _0331_ VGND controller.inst_mem.mem_data\[153\] net586 sg13g2_o21ai_1
Xhold1 controller.inst_mem.mem_data\[64\] VPWR VGND net328 sg13g2_dlygate4sd3_1
X_3248__182 VPWR VGND net182 sg13g2_tiehi
X_2875_ net641 VPWR _0929_ VGND controller.const_data\[30\] net576 sg13g2_o21ai_1
X_1826_ VPWR _1177_ net839 VGND sg13g2_inv_1
Xhold401 controller.alu_buffer.buffer\[20\] VPWR VGND net948 sg13g2_dlygate4sd3_1
X_2944_ VGND VPWR _0997_ net549 _0272_ _0963_ sg13g2_a21oi_1
X_3023__78 VPWR VGND net78 sg13g2_tiehi
X_1688_ VPWR _1039_ net718 VGND sg13g2_inv_1
Xhold434 _0154_ VPWR VGND net981 sg13g2_dlygate4sd3_1
Xhold423 _0161_ VPWR VGND net970 sg13g2_dlygate4sd3_1
Xhold412 _0166_ VPWR VGND net959 sg13g2_dlygate4sd3_1
X_1757_ VPWR _1108_ net438 VGND sg13g2_inv_1
X_3075__263 VPWR VGND net263 sg13g2_tiehi
X_2309_ _0451_ _0452_ _0453_ _0454_ _0455_ VPWR VGND sg13g2_nor4_1
X_2660_ net540 VPWR _0776_ VGND net947 net444 sg13g2_o21ai_1
X_3212_ net322 VGND VPWR _0235_ controller.const_data\[27\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2591_ _0711_ _1064_ net455 VPWR VGND sg13g2_nand2_1
XFILLER_4_481 VPWR VGND sg13g2_fill_1
X_3143_ net85 VGND VPWR net959 controller.alu_buffer.buffer\[17\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
X_2025_ net625 VPWR _1339_ VGND net828 net550 sg13g2_o21ai_1
X_3074_ net265 VGND VPWR net698 controller.inst_mem.mem_data\[178\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_35_385 VPWR VGND sg13g2_fill_2
X_2927_ net648 VPWR _0955_ VGND net804 net593 sg13g2_o21ai_1
X_2858_ VGND VPWR _1040_ net614 _0229_ _0920_ sg13g2_a21oi_1
X_2789_ VGND VPWR net396 net451 _0878_ _0877_ sg13g2_a21oi_1
X_1809_ VPWR _1160_ net435 VGND sg13g2_inv_1
Xhold231 controller.inst_mem.mem_data\[83\] VPWR VGND net778 sg13g2_dlygate4sd3_1
Xhold242 controller.inst_mem.mem_data\[87\] VPWR VGND net789 sg13g2_dlygate4sd3_1
Xhold253 controller.inst_mem.mem_data\[34\] VPWR VGND net800 sg13g2_dlygate4sd3_1
Xhold220 controller.inst_mem.mem_data\[67\] VPWR VGND net767 sg13g2_dlygate4sd3_1
Xhold286 _0211_ VPWR VGND net833 sg13g2_dlygate4sd3_1
Xhold275 controller.const_data\[28\] VPWR VGND net822 sg13g2_dlygate4sd3_1
Xhold264 controller.const_data\[24\] VPWR VGND net811 sg13g2_dlygate4sd3_1
Xhold297 controller.extended_jump_target\[0\] VPWR VGND net844 sg13g2_dlygate4sd3_1
XFILLER_5_267 VPWR VGND sg13g2_fill_2
XFILLER_5_278 VPWR VGND sg13g2_fill_1
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_32_355 VPWR VGND sg13g2_fill_1
X_2712_ VGND VPWR net445 _0815_ _0187_ _0816_ sg13g2_a21oi_1
X_2574_ _0696_ net960 _1297_ VPWR VGND sg13g2_xnor2_1
X_2643_ net519 controller.inst_mem.mem_data\[140\] net515 _0759_ VPWR VGND sg13g2_a21o_1
X_3126_ net153 VGND VPWR net968 controller.alu_buffer.buffer\[8\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_2008_ VGND VPWR _1196_ net600 _0020_ _1330_ sg13g2_a21oi_1
X_3057_ net299 VGND VPWR _0080_ controller.inst_mem.mem_data\[161\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
Xfanout541 net542 net541 VPWR VGND sg13g2_buf_8
Xfanout530 net983 net530 VPWR VGND sg13g2_buf_8
Xfanout574 net579 net574 VPWR VGND sg13g2_buf_8
Xfanout585 net586 net585 VPWR VGND sg13g2_buf_8
Xfanout552 net553 net552 VPWR VGND sg13g2_buf_2
Xfanout596 net597 net596 VPWR VGND sg13g2_buf_8
Xfanout563 net564 net563 VPWR VGND sg13g2_buf_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_14_388 VPWR VGND sg13g2_fill_1
X_2290_ _1087_ _0430_ _0436_ VPWR VGND sg13g2_nor2_1
XFILLER_49_296 VPWR VGND sg13g2_fill_1
XFILLER_45_491 VPWR VGND sg13g2_decap_8
XFILLER_37_447 VPWR VGND sg13g2_decap_8
X_2626_ _0742_ net496 controller.inst_mem.mem_data\[94\] net512 controller.inst_mem.mem_data\[166\]
+ VPWR VGND sg13g2_a22oi_1
X_2557_ VPWR VGND net466 net461 _0681_ net945 _0682_ net481 sg13g2_a221oi_1
X_2488_ VGND VPWR _0621_ _0624_ _0154_ _0625_ sg13g2_a21oi_1
X_3109_ net195 VGND VPWR _0132_ controller.extended_then_action\[1\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
X_3194__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_36_82 VPWR VGND sg13g2_fill_2
XFILLER_34_406 VPWR VGND sg13g2_fill_1
Xinput13 uio_in[6] net13 VPWR VGND sg13g2_buf_1
X_1790_ VPWR _1141_ net703 VGND sg13g2_inv_1
X_2411_ _0554_ controller.inst_mem.mem_data\[121\] net499 VPWR VGND sg13g2_nand2_1
X_2273_ _0419_ _0418_ controller.counter2.counter_0\[15\] VPWR VGND sg13g2_nand2b_1
X_2342_ _0488_ controller.inst_mem.mem_data\[179\] net502 VPWR VGND sg13g2_nand2_1
XFILLER_33_472 VPWR VGND sg13g2_decap_8
X_1988_ VGND VPWR _1206_ net566 _0010_ _1320_ sg13g2_a21oi_1
XFILLER_20_144 VPWR VGND sg13g2_fill_1
X_2609_ _0725_ _0479_ controller.inst_mem.mem_data\[141\] net513 controller.inst_mem.mem_data\[165\]
+ VPWR VGND sg13g2_a22oi_1
X_3085__243 VPWR VGND net243 sg13g2_tiehi
XFILLER_0_0 VPWR VGND sg13g2_fill_2
X_2960_ VGND VPWR _0989_ net617 _0280_ _0971_ sg13g2_a21oi_1
X_1842_ VPWR _1193_ net868 VGND sg13g2_inv_1
X_1773_ VPWR _1124_ net825 VGND sg13g2_inv_1
X_2891_ net631 VPWR _0937_ VGND controller.inst_mem.mem_data\[38\] net558 sg13g2_o21ai_1
X_3035__54 VPWR VGND net54 sg13g2_tiehi
X_1911_ VGND VPWR controller.output_controller.keep\[0\] _1261_ _1262_ _1249_ sg13g2_a21oi_1
X_2187_ net656 VPWR _0369_ VGND controller.inst_mem.mem_data\[191\] net610 sg13g2_o21ai_1
X_2325_ _0471_ net2 _0448_ VPWR VGND sg13g2_nand2b_1
X_2256_ VGND VPWR _1072_ net589 _0144_ _0403_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_32 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_3_162 VPWR VGND sg13g2_fill_1
XFILLER_3_151 VPWR VGND sg13g2_fill_1
X_2041_ net655 VPWR _0296_ VGND net768 net606 sg13g2_o21ai_1
X_3090_ net233 VGND VPWR _0113_ controller.inst_mem.mem_data\[194\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_2110_ VGND VPWR _1145_ net592 _0071_ _0330_ sg13g2_a21oi_1
Xhold2 _0273_ VPWR VGND net329 sg13g2_dlygate4sd3_1
XFILLER_47_394 VPWR VGND sg13g2_decap_8
X_2943_ net625 VPWR _0963_ VGND net328 net549 sg13g2_o21ai_1
X_2874_ VGND VPWR _1032_ net576 _0237_ _0928_ sg13g2_a21oi_1
Xhold435 controller.alu_buffer.buffer\[6\] VPWR VGND net982 sg13g2_dlygate4sd3_1
Xhold424 controller.alu_buffer.buffer\[0\] VPWR VGND net971 sg13g2_dlygate4sd3_1
X_1825_ VPWR _1176_ net760 VGND sg13g2_inv_1
X_1756_ VPWR _1107_ net717 VGND sg13g2_inv_1
Xhold413 controller.alu_buffer.buffer\[21\] VPWR VGND net960 sg13g2_dlygate4sd3_1
Xhold402 _0169_ VPWR VGND net949 sg13g2_dlygate4sd3_1
X_1687_ VPWR _1038_ net840 VGND sg13g2_inv_1
X_2308_ _1109_ _1223_ _0454_ VPWR VGND sg13g2_nor2_1
X_2239_ net660 VPWR _0395_ VGND net878 net616 sg13g2_o21ai_1
XFILLER_44_375 VPWR VGND sg13g2_fill_1
X_2590_ net456 _0708_ _0709_ _0710_ VPWR VGND sg13g2_or3_1
X_3211_ net41 VGND VPWR net688 controller.const_data\[26\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_3142_ net89 VGND VPWR net966 controller.alu_buffer.buffer\[16\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
XFILLER_39_169 VPWR VGND sg13g2_fill_2
X_3111__191 VPWR VGND net191 sg13g2_tiehi
X_3073_ net267 VGND VPWR _0096_ controller.inst_mem.mem_data\[177\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
X_2024_ VGND VPWR _1188_ net555 _0028_ _1338_ sg13g2_a21oi_1
X_2857_ net658 VPWR _0920_ VGND net718 net612 sg13g2_o21ai_1
X_2926_ VGND VPWR _1006_ net589 _0263_ _0954_ sg13g2_a21oi_1
X_2788_ VGND VPWR _1277_ _0876_ _0877_ net451 sg13g2_a21oi_1
Xhold221 controller.inst_mem.mem_data\[118\] VPWR VGND net768 sg13g2_dlygate4sd3_1
Xhold254 controller.inst_mem.mem_data\[94\] VPWR VGND net801 sg13g2_dlygate4sd3_1
Xhold232 controller.inst_mem.mem_data\[117\] VPWR VGND net779 sg13g2_dlygate4sd3_1
Xhold276 controller.inst_mem.mem_data\[154\] VPWR VGND net823 sg13g2_dlygate4sd3_1
X_1739_ VPWR _1090_ net701 VGND sg13g2_inv_1
X_1808_ VPWR _1159_ net351 VGND sg13g2_inv_1
Xhold210 controller.inst_mem.mem_data\[112\] VPWR VGND net757 sg13g2_dlygate4sd3_1
Xhold265 controller.inst_mem.mem_data\[53\] VPWR VGND net812 sg13g2_dlygate4sd3_1
Xhold287 controller.inst_mem.mem_data\[187\] VPWR VGND net834 sg13g2_dlygate4sd3_1
Xhold243 controller.inst_mem.mem_data\[195\] VPWR VGND net790 sg13g2_dlygate4sd3_1
XFILLER_45_117 VPWR VGND sg13g2_fill_1
Xhold298 _0120_ VPWR VGND net845 sg13g2_dlygate4sd3_1
XFILLER_26_331 VPWR VGND sg13g2_fill_2
X_3212__322 VPWR VGND net322 sg13g2_tiehi
XFILLER_49_445 VPWR VGND sg13g2_decap_8
X_3169__276 VPWR VGND net276 sg13g2_tiehi
X_2711_ net541 VPWR _0816_ VGND net897 net445 sg13g2_o21ai_1
X_2642_ _0758_ _1016_ net516 VPWR VGND sg13g2_nand2_1
X_2573_ controller.alu_buffer.buffer\[21\] _1297_ _0695_ VPWR VGND sg13g2_nor2_1
X_3125_ net157 VGND VPWR net987 controller.inst_mem.addr\[2\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3224__226 VPWR VGND net226 sg13g2_tiehi
X_2007_ net652 VPWR _1330_ VGND controller.inst_mem.mem_data\[101\] net600 sg13g2_o21ai_1
X_3044__325 VPWR VGND net325 sg13g2_tiehi
X_3056_ net301 VGND VPWR _0079_ controller.inst_mem.mem_data\[160\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_2909_ net657 VPWR _0946_ VGND net413 net606 sg13g2_o21ai_1
Xfanout542 _0502_ net542 VPWR VGND sg13g2_buf_8
Xfanout531 net532 net531 VPWR VGND sg13g2_buf_8
Xfanout520 net522 net520 VPWR VGND sg13g2_buf_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
Xfanout575 net579 net575 VPWR VGND sg13g2_buf_8
Xfanout586 net587 net586 VPWR VGND sg13g2_buf_8
Xfanout597 net605 net597 VPWR VGND sg13g2_buf_8
Xfanout553 net554 net553 VPWR VGND sg13g2_buf_2
Xfanout564 net567 net564 VPWR VGND sg13g2_buf_8
X_3125__157 VPWR VGND net157 sg13g2_tiehi
X_3095__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_45_470 VPWR VGND sg13g2_decap_8
X_2487_ net539 VPWR _0625_ VGND net528 net460 sg13g2_o21ai_1
X_2625_ net521 controller.inst_mem.mem_data\[142\] _1231_ _0741_ VPWR VGND sg13g2_a21o_1
X_2556_ _0676_ net952 _0681_ VPWR VGND sg13g2_xor2_1
X_3108_ net197 VGND VPWR _0131_ controller.extended_then_action\[0\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_43_429 VPWR VGND sg13g2_decap_8
X_3039_ net46 VGND VPWR net369 controller.inst_mem.mem_data\[143\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_7_308 VPWR VGND sg13g2_fill_1
Xinput14 uio_in[7] net14 VPWR VGND sg13g2_buf_1
XFILLER_42_484 VPWR VGND sg13g2_decap_8
X_2410_ VGND VPWR _0439_ _0552_ _0553_ _0475_ sg13g2_a21oi_1
X_2341_ _0487_ net523 controller.inst_mem.extended_word\[3\] net506 controller.inst_mem.mem_data\[59\]
+ VPWR VGND sg13g2_a22oi_1
X_2272_ net893 net897 _0414_ _0416_ _0418_ VPWR VGND sg13g2_nor4_1
XFILLER_37_289 VPWR VGND sg13g2_fill_1
X_1987_ net633 VPWR _1320_ VGND controller.inst_mem.mem_data\[91\] net566 sg13g2_o21ai_1
X_2539_ _0667_ _0666_ net466 net456 controller.alu_buffer.buffer\[7\] VPWR VGND sg13g2_a22oi_1
X_2608_ _0724_ net526 controller.extended_then_action\[1\] net509 controller.inst_mem.mem_data\[69\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_3_355 VPWR VGND sg13g2_fill_1
X_2890_ VGND VPWR _1024_ net561 _0245_ _0936_ sg13g2_a21oi_1
X_1910_ _1235_ _1242_ _1261_ VPWR VGND sg13g2_nor2b_1
X_1772_ VPWR _1123_ net810 VGND sg13g2_inv_1
X_1841_ VPWR _1192_ net388 VGND sg13g2_inv_1
XFILLER_8_32 VPWR VGND sg13g2_fill_1
X_2324_ _1280_ _1300_ _0448_ _0470_ VPWR VGND sg13g2_mux2_1
XFILLER_26_0 VPWR VGND sg13g2_fill_2
X_2186_ VGND VPWR _1107_ net606 _0109_ _0368_ sg13g2_a21oi_1
X_2255_ net647 VPWR _0403_ VGND controller.extended_state\[1\] net589 sg13g2_o21ai_1
X_3121__171 VPWR VGND net171 sg13g2_tiehi
Xheichips25_can_lehmann_fsm_33 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_0_303 VPWR VGND sg13g2_fill_2
X_3232__155 VPWR VGND net155 sg13g2_tiehi
X_3243__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_47_373 VPWR VGND sg13g2_decap_8
Xhold3 controller.inst_mem.mem_data\[141\] VPWR VGND net330 sg13g2_dlygate4sd3_1
X_2040_ VGND VPWR _1180_ net573 _0036_ _0295_ sg13g2_a21oi_1
X_2873_ net641 VPWR _0928_ VGND net440 net576 sg13g2_o21ai_1
X_2942_ VGND VPWR _0998_ net548 _0271_ _0962_ sg13g2_a21oi_1
X_1686_ VPWR _1037_ net820 VGND sg13g2_inv_1
Xhold414 controller.alu_buffer.buffer\[4\] VPWR VGND net961 sg13g2_dlygate4sd3_1
Xhold436 controller.alu_buffer.buffer\[1\] VPWR VGND net983 sg13g2_dlygate4sd3_1
Xhold425 _0150_ VPWR VGND net972 sg13g2_dlygate4sd3_1
X_1824_ VPWR _1175_ net737 VGND sg13g2_inv_1
X_1755_ VPWR _1106_ net380 VGND sg13g2_inv_1
Xhold403 controller.alu_buffer.buffer\[14\] VPWR VGND net950 sg13g2_dlygate4sd3_1
X_2238_ VGND VPWR _1081_ net611 _0135_ _0394_ sg13g2_a21oi_1
X_2307_ net531 _1181_ _1225_ _0453_ VPWR VGND sg13g2_nor3_1
X_3227__202 VPWR VGND net202 sg13g2_tiehi
X_2169_ net625 VPWR _0360_ VGND controller.inst_mem.mem_data\[182\] net548 sg13g2_o21ai_1
XFILLER_21_251 VPWR VGND sg13g2_fill_1
XFILLER_21_284 VPWR VGND sg13g2_fill_2
X_3054__305 VPWR VGND net305 sg13g2_tiehi
X_3022__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_44_354 VPWR VGND sg13g2_fill_2
XFILLER_8_233 VPWR VGND sg13g2_fill_2
XFILLER_12_295 VPWR VGND sg13g2_fill_2
X_3210_ net49 VGND VPWR _0233_ controller.const_data\[25\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3141_ net93 VGND VPWR net923 controller.alu_buffer.buffer\[15\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_2023_ net628 VPWR _1338_ VGND net855 net555 sg13g2_o21ai_1
X_3072_ net269 VGND VPWR net700 controller.inst_mem.mem_data\[176\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_2856_ VGND VPWR _1041_ net612 _0228_ _0919_ sg13g2_a21oi_1
X_2925_ net653 VPWR _0954_ VGND controller.inst_mem.mem_data\[55\] net598 sg13g2_o21ai_1
X_1807_ VPWR _1158_ net355 VGND sg13g2_inv_1
Xhold277 controller.const_data\[7\] VPWR VGND net824 sg13g2_dlygate4sd3_1
X_2787_ _0876_ net883 _1275_ VPWR VGND sg13g2_nand2_1
Xhold222 _0038_ VPWR VGND net769 sg13g2_dlygate4sd3_1
X_1738_ VPWR _1089_ net782 VGND sg13g2_inv_1
Xhold266 controller.inst_mem.mem_data\[192\] VPWR VGND net813 sg13g2_dlygate4sd3_1
Xhold255 _0014_ VPWR VGND net802 sg13g2_dlygate4sd3_1
X_1669_ VPWR _1020_ net722 VGND sg13g2_inv_1
Xhold233 controller.inst_mem.mem_data\[170\] VPWR VGND net780 sg13g2_dlygate4sd3_1
Xhold211 controller.inst_mem.mem_data\[62\] VPWR VGND net758 sg13g2_dlygate4sd3_1
Xhold299 controller.inst_mem.mem_data\[184\] VPWR VGND net846 sg13g2_dlygate4sd3_1
Xhold288 controller.inst_mem.mem_data\[76\] VPWR VGND net835 sg13g2_dlygate4sd3_1
Xhold200 controller.inst_mem.mem_data\[140\] VPWR VGND net747 sg13g2_dlygate4sd3_1
Xhold244 _0115_ VPWR VGND net791 sg13g2_dlygate4sd3_1
X_2986__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_41_357 VPWR VGND sg13g2_fill_2
XFILLER_49_424 VPWR VGND sg13g2_decap_8
X_3176__248 VPWR VGND net248 sg13g2_tiehi
X_2710_ _0815_ net449 _0814_ _0767_ net681 VPWR VGND sg13g2_a22oi_1
X_2572_ VPWR VGND net956 net461 net481 net948 _0694_ net470 sg13g2_a221oi_1
X_2641_ _0755_ _0756_ net487 _0757_ VPWR VGND sg13g2_nand3_1
X_3055_ net303 VGND VPWR net795 controller.inst_mem.mem_data\[159\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_3124_ net161 VGND VPWR net979 controller.inst_mem.addr\[1\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_2006_ VGND VPWR _1197_ net601 _0019_ _1329_ sg13g2_a21oi_1
X_2839_ net640 VPWR _0911_ VGND net372 net577 sg13g2_o21ai_1
X_2908_ VGND VPWR _1015_ net574 _0254_ _0945_ sg13g2_a21oi_1
Xfanout543 net545 net543 VPWR VGND sg13g2_buf_8
Xfanout554 net568 net554 VPWR VGND sg13g2_buf_8
Xfanout521 net522 net521 VPWR VGND sg13g2_buf_1
Xfanout532 net986 net532 VPWR VGND sg13g2_buf_8
Xfanout565 net567 net565 VPWR VGND sg13g2_buf_8
Xfanout510 net513 net510 VPWR VGND sg13g2_buf_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
Xfanout576 net578 net576 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_38_clk clknet_3_0__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
Xfanout587 net591 net587 VPWR VGND sg13g2_buf_8
Xfanout598 net604 net598 VPWR VGND sg13g2_buf_8
X_3132__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_1_272 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_29_clk clknet_3_4__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_17_140 VPWR VGND sg13g2_fill_2
X_2624_ _0740_ net500 controller.inst_mem.mem_data\[118\] net508 controller.inst_mem.mem_data\[70\]
+ VPWR VGND sg13g2_a22oi_1
X_2486_ _0624_ _0623_ net468 net457 net11 VPWR VGND sg13g2_a22oi_1
X_2555_ controller.alu_buffer.buffer\[18\] _0676_ _0680_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_408 VPWR VGND sg13g2_decap_8
X_3107_ net199 VGND VPWR _0130_ controller.extended_cond.opcode\[2\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_3038_ net48 VGND VPWR net331 controller.inst_mem.mem_data\[142\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_36_482 VPWR VGND sg13g2_decap_8
XFILLER_23_110 VPWR VGND sg13g2_fill_1
XFILLER_42_463 VPWR VGND sg13g2_decap_8
XFILLER_10_382 VPWR VGND sg13g2_fill_2
X_3062__289 VPWR VGND net289 sg13g2_tiehi
X_2271_ _0415_ _0416_ _0417_ VPWR VGND sg13g2_nor2_1
X_2340_ net515 _1024_ _0484_ _0486_ VPWR VGND sg13g2_a21o_2
X_3108__197 VPWR VGND net197 sg13g2_tiehi
X_1986_ VGND VPWR _1207_ net564 _0009_ _1319_ sg13g2_a21oi_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_2607_ _0723_ net497 controller.inst_mem.mem_data\[93\] net501 controller.inst_mem.mem_data\[117\]
+ VPWR VGND sg13g2_a22oi_1
X_2469_ net539 VPWR _0610_ VGND net530 net460 sg13g2_o21ai_1
X_2538_ _1294_ VPWR _0666_ VGND _1064_ _0660_ sg13g2_o21ai_1
XFILLER_34_216 VPWR VGND sg13g2_fill_2
X_1840_ VPWR _1191_ net805 VGND sg13g2_inv_1
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_30_477 VPWR VGND sg13g2_fill_2
X_1771_ VPWR _1122_ net738 VGND sg13g2_inv_1
XFILLER_38_500 VPWR VGND sg13g2_decap_8
X_2323_ VPWR VGND _0468_ _0465_ _0467_ _0419_ _0469_ _0458_ sg13g2_a221oi_1
X_2254_ VGND VPWR _1073_ net589 _0143_ _0402_ sg13g2_a21oi_1
X_2185_ net655 VPWR _0368_ VGND net380 net606 sg13g2_o21ai_1
XFILLER_19_0 VPWR VGND sg13g2_fill_2
X_1969_ net643 VPWR _1311_ VGND net677 net586 sg13g2_o21ai_1
Xheichips25_can_lehmann_fsm_23 VPWR VGND uio_oe[0] sg13g2_tielo
Xheichips25_can_lehmann_fsm_34 VPWR VGND uio_out[3] sg13g2_tielo
X_2996__132 VPWR VGND net132 sg13g2_tiehi
Xhold4 _0061_ VPWR VGND net331 sg13g2_dlygate4sd3_1
XFILLER_35_503 VPWR VGND sg13g2_decap_4
X_2872_ VGND VPWR _1033_ net612 _0236_ _0927_ sg13g2_a21oi_1
X_1823_ VPWR _1174_ net362 VGND sg13g2_inv_1
X_2941_ net625 VPWR _0962_ VGND controller.inst_mem.mem_data\[63\] net546 sg13g2_o21ai_1
XFILLER_22_219 VPWR VGND sg13g2_fill_1
X_3190__192 VPWR VGND net192 sg13g2_tiehi
Xhold415 _0155_ VPWR VGND net962 sg13g2_dlygate4sd3_1
Xhold437 controller.alu_buffer.buffer\[0\] VPWR VGND net984 sg13g2_dlygate4sd3_1
Xhold426 controller.alu_buffer.buffer\[7\] VPWR VGND net973 sg13g2_dlygate4sd3_1
X_1685_ VPWR _1036_ net811 VGND sg13g2_inv_1
X_1754_ VPWR _1105_ net394 VGND sg13g2_inv_1
Xhold404 _0163_ VPWR VGND net951 sg13g2_dlygate4sd3_1
X_2237_ net656 VPWR _0394_ VGND net881 net611 sg13g2_o21ai_1
X_2306_ net519 controller.inst_mem.mem_data\[139\] net515 _0452_ VPWR VGND sg13g2_a21o_1
XFILLER_41_506 VPWR VGND sg13g2_fill_2
XFILLER_38_385 VPWR VGND sg13g2_fill_1
X_2168_ VGND VPWR _1116_ net555 _0100_ _0359_ sg13g2_a21oi_1
X_2099_ net653 VPWR _0325_ VGND net436 net598 sg13g2_o21ai_1
X_3128__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_44_366 VPWR VGND sg13g2_fill_2
XFILLER_32_506 VPWR VGND sg13g2_fill_2
X_3140_ net97 VGND VPWR net951 controller.alu_buffer.buffer\[14\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_3071_ net271 VGND VPWR _0094_ controller.inst_mem.mem_data\[175\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_2022_ VGND VPWR _1189_ net559 _0027_ _1337_ sg13g2_a21oi_1
X_2855_ net658 VPWR _0919_ VGND controller.const_data\[20\] net612 sg13g2_o21ai_1
X_2786_ VGND VPWR net478 _0874_ _0202_ _0875_ sg13g2_a21oi_1
Xhold201 controller.inst_mem.mem_data\[35\] VPWR VGND net748 sg13g2_dlygate4sd3_1
X_2924_ VGND VPWR _1007_ net589 _0262_ _0953_ sg13g2_a21oi_1
X_1806_ VPWR _1157_ net411 VGND sg13g2_inv_1
Xhold256 controller.inst_mem.mem_data\[70\] VPWR VGND net803 sg13g2_dlygate4sd3_1
X_1737_ VPWR _1088_ net761 VGND sg13g2_inv_1
X_1668_ VPWR _1019_ net856 VGND sg13g2_inv_1
Xhold212 _0271_ VPWR VGND net759 sg13g2_dlygate4sd3_1
Xhold223 controller.inst_mem.mem_data\[89\] VPWR VGND net770 sg13g2_dlygate4sd3_1
Xhold278 controller.inst_mem.mem_data\[172\] VPWR VGND net825 sg13g2_dlygate4sd3_1
Xhold267 controller.inst_mem.mem_data\[186\] VPWR VGND net814 sg13g2_dlygate4sd3_1
Xhold245 controller.inst_mem.mem_data\[75\] VPWR VGND net792 sg13g2_dlygate4sd3_1
Xhold289 controller.inst_mem.mem_data\[100\] VPWR VGND net836 sg13g2_dlygate4sd3_1
Xhold234 controller.inst_mem.mem_data\[143\] VPWR VGND net781 sg13g2_dlygate4sd3_1
XFILLER_49_403 VPWR VGND sg13g2_decap_8
X_2640_ controller.extended_then_action\[0\] net490 net489 _0756_ VPWR VGND sg13g2_or3_1
X_2571_ VGND VPWR _0690_ _0692_ _0169_ _0693_ sg13g2_a21oi_1
X_3072__269 VPWR VGND net269 sg13g2_tiehi
XFILLER_48_491 VPWR VGND sg13g2_decap_8
X_3054_ net305 VGND VPWR _0077_ controller.inst_mem.mem_data\[158\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_3123_ net165 VGND VPWR _0146_ controller.inst_mem.addr\[0\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_2005_ net651 VPWR _1329_ VGND controller.inst_mem.mem_data\[100\] net601 sg13g2_o21ai_1
X_2907_ net639 VPWR _0945_ VGND controller.inst_mem.mem_data\[46\] net574 sg13g2_o21ai_1
XFILLER_23_347 VPWR VGND sg13g2_fill_1
X_2838_ VGND VPWR _1050_ net571 _0219_ _0910_ sg13g2_a21oi_1
X_2769_ net543 VPWR _0862_ VGND net932 net476 sg13g2_o21ai_1
XFILLER_46_406 VPWR VGND sg13g2_decap_8
Xfanout577 net579 net577 VPWR VGND sg13g2_buf_8
Xfanout544 net545 net544 VPWR VGND sg13g2_buf_8
Xfanout555 net557 net555 VPWR VGND sg13g2_buf_8
X_3118__177 VPWR VGND net177 sg13g2_tiehi
Xfanout533 net978 net533 VPWR VGND sg13g2_buf_8
Xfanout588 net589 net588 VPWR VGND sg13g2_buf_8
Xfanout566 net567 net566 VPWR VGND sg13g2_buf_8
Xfanout511 net513 net511 VPWR VGND sg13g2_buf_8
Xfanout522 _1230_ net522 VPWR VGND sg13g2_buf_2
Xfanout599 net603 net599 VPWR VGND sg13g2_buf_8
Xfanout500 net501 net500 VPWR VGND sg13g2_buf_8
XFILLER_39_480 VPWR VGND sg13g2_decap_8
X_3216__290 VPWR VGND net290 sg13g2_tiehi
X_2623_ controller.extended_then_action\[2\] _0738_ net488 _0739_ VPWR VGND sg13g2_mux2_1
X_2554_ VGND VPWR _0675_ _0678_ _0166_ _0679_ sg13g2_a21oi_1
X_2485_ _1283_ net528 _0623_ VPWR VGND sg13g2_xor2_1
XFILLER_36_461 VPWR VGND sg13g2_decap_8
X_3106_ net201 VGND VPWR net937 controller.extended_cond.opcode\[1\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_3228__194 VPWR VGND net194 sg13g2_tiehi
X_3037_ net50 VGND VPWR _0060_ controller.inst_mem.mem_data\[141\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_11_306 VPWR VGND sg13g2_fill_1
XFILLER_42_442 VPWR VGND sg13g2_decap_8
X_2270_ VGND VPWR _0416_ controller.counter2.counter_0\[12\] controller.counter2.counter_0\[13\]
+ sg13g2_or2_1
XFILLER_37_225 VPWR VGND sg13g2_fill_2
XFILLER_33_486 VPWR VGND sg13g2_decap_8
X_1985_ net633 VPWR _1319_ VGND net423 net562 sg13g2_o21ai_1
X_2606_ _0722_ net487 _0720_ _0721_ VPWR VGND sg13g2_and3_1
X_2537_ VPWR VGND controller.alu_buffer.buffer\[16\] net461 net481 controller.alu_buffer.buffer\[14\]
+ _0665_ net470 sg13g2_a221oi_1
X_2468_ VPWR VGND net529 net463 net483 net971 _0609_ net473 sg13g2_a221oi_1
X_2399_ _0539_ _0540_ _0538_ _0542_ VPWR VGND _0541_ sg13g2_nand4_1
X_3165__292 VPWR VGND net292 sg13g2_tiehi
XFILLER_28_258 VPWR VGND sg13g2_fill_1
XFILLER_24_475 VPWR VGND sg13g2_fill_2
XFILLER_47_73 VPWR VGND sg13g2_fill_1
X_1770_ VPWR _1121_ net699 VGND sg13g2_inv_1
XFILLER_8_78 VPWR VGND sg13g2_fill_2
X_2322_ VGND VPWR net3 _0448_ _0468_ _0457_ sg13g2_a21oi_1
X_2253_ net647 VPWR _0402_ VGND net376 net589 sg13g2_o21ai_1
X_2184_ VGND VPWR _1108_ net573 _0108_ _0367_ sg13g2_a21oi_1
X_1899_ VPWR VGND controller.inst_mem.mem_data\[134\] net514 net519 controller.inst_mem.mem_data\[86\]
+ _1250_ net494 sg13g2_a221oi_1
X_1968_ VGND VPWR _0980_ net586 _0000_ _1310_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_24 VPWR VGND uio_oe[1] sg13g2_tielo
Xheichips25_can_lehmann_fsm_35 VPWR VGND uio_out[4] sg13g2_tielo
X_3100__213 VPWR VGND net213 sg13g2_tiehi
Xhold5 controller.inst_mem.mem_data\[144\] VPWR VGND net332 sg13g2_dlygate4sd3_1
X_2940_ VGND VPWR _0999_ net553 _0270_ _0961_ sg13g2_a21oi_1
X_3179__236 VPWR VGND net236 sg13g2_tiehi
X_2871_ net658 VPWR _0927_ VGND controller.const_data\[28\] net612 sg13g2_o21ai_1
X_1753_ VPWR _1104_ net813 VGND sg13g2_inv_1
X_3001__122 VPWR VGND net122 sg13g2_tiehi
X_1822_ VPWR _1173_ net742 VGND sg13g2_inv_1
X_1684_ VPWR _1035_ net687 VGND sg13g2_inv_1
Xhold427 _0157_ VPWR VGND net974 sg13g2_dlygate4sd3_1
Xhold416 controller.alu_buffer.buffer\[9\] VPWR VGND net963 sg13g2_dlygate4sd3_1
XFILLER_31_0 VPWR VGND sg13g2_fill_2
Xhold438 controller.inst_mem.addr\[0\] VPWR VGND net985 sg13g2_dlygate4sd3_1
Xhold405 controller.alu_buffer.buffer\[18\] VPWR VGND net952 sg13g2_dlygate4sd3_1
XFILLER_38_375 VPWR VGND sg13g2_fill_1
X_2236_ VGND VPWR _1082_ net608 _0134_ _0393_ sg13g2_a21oi_1
X_2167_ net629 VPWR _0359_ VGND controller.inst_mem.mem_data\[181\] net555 sg13g2_o21ai_1
X_2305_ net531 _1205_ _1221_ _0451_ VPWR VGND sg13g2_nor3_1
X_2098_ VGND VPWR _1151_ net615 _0065_ _0324_ sg13g2_a21oi_1
X_3082__249 VPWR VGND net249 sg13g2_tiehi
XFILLER_28_31 VPWR VGND sg13g2_fill_1
XFILLER_44_356 VPWR VGND sg13g2_fill_1
XFILLER_12_286 VPWR VGND sg13g2_fill_1
X_3135__117 VPWR VGND net117 sg13g2_tiehi
XFILLER_4_474 VPWR VGND sg13g2_fill_2
X_2021_ net630 VPWR _1337_ VGND controller.inst_mem.mem_data\[108\] net559 sg13g2_o21ai_1
X_3070_ net273 VGND VPWR _0093_ controller.inst_mem.mem_data\[174\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_23_507 VPWR VGND sg13g2_fill_1
X_2923_ net647 VPWR _0953_ VGND net726 net589 sg13g2_o21ai_1
X_2854_ VGND VPWR _1042_ net576 _0227_ _0918_ sg13g2_a21oi_1
X_2785_ net543 VPWR _0875_ VGND net907 net478 sg13g2_o21ai_1
Xhold213 controller.inst_mem.mem_data\[120\] VPWR VGND net760 sg13g2_dlygate4sd3_1
X_1736_ VPWR _1087_ net936 VGND sg13g2_inv_1
Xhold224 controller.inst_mem.mem_data\[152\] VPWR VGND net771 sg13g2_dlygate4sd3_1
Xhold235 controller.inst_mem.extended_word\[7\] VPWR VGND net782 sg13g2_dlygate4sd3_1
Xhold202 _0244_ VPWR VGND net749 sg13g2_dlygate4sd3_1
X_1805_ VPWR _1156_ net747 VGND sg13g2_inv_1
X_1667_ VPWR _1018_ net740 VGND sg13g2_inv_1
Xhold257 controller.inst_mem.mem_data\[56\] VPWR VGND net804 sg13g2_dlygate4sd3_1
Xhold246 _0284_ VPWR VGND net793 sg13g2_dlygate4sd3_1
Xhold279 controller.inst_mem.mem_data\[77\] VPWR VGND net826 sg13g2_dlygate4sd3_1
Xhold268 _0106_ VPWR VGND net815 sg13g2_dlygate4sd3_1
X_3199_ net143 VGND VPWR _0222_ controller.const_data\[14\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2219_ net626 VPWR _0385_ VGND controller.inst_mem.extended_word\[7\] net549 sg13g2_o21ai_1
XFILLER_14_507 VPWR VGND sg13g2_fill_1
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_17_345 VPWR VGND sg13g2_fill_2
X_2570_ net537 VPWR _0693_ VGND net948 net458 sg13g2_o21ai_1
X_3122_ net169 VGND VPWR net752 controller.extended_state\[2\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_48_470 VPWR VGND sg13g2_decap_8
X_2004_ VGND VPWR _1198_ net620 _0018_ _1328_ sg13g2_a21oi_1
X_3053_ net307 VGND VPWR _0076_ controller.inst_mem.mem_data\[157\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_2906_ VGND VPWR _1016_ net574 _0253_ _0944_ sg13g2_a21oi_1
X_2837_ net640 VPWR _0910_ VGND net681 net571 sg13g2_o21ai_1
X_2699_ VGND VPWR net445 _0805_ _0184_ _0806_ sg13g2_a21oi_1
X_2768_ VGND VPWR net820 net452 _0861_ _0860_ sg13g2_a21oi_1
X_1719_ VPWR _1070_ net535 VGND sg13g2_inv_1
Xfanout578 net579 net578 VPWR VGND sg13g2_buf_1
Xfanout545 _0502_ net545 VPWR VGND sg13g2_buf_8
Xfanout556 net557 net556 VPWR VGND sg13g2_buf_1
Xfanout589 net591 net589 VPWR VGND sg13g2_buf_8
Xfanout534 controller.inst_mem.addr\[1\] net534 VPWR VGND sg13g2_buf_8
Xfanout567 net568 net567 VPWR VGND sg13g2_buf_8
Xfanout501 _1226_ net501 VPWR VGND sg13g2_buf_8
Xfanout523 net526 net523 VPWR VGND sg13g2_buf_8
Xfanout512 net513 net512 VPWR VGND sg13g2_buf_2
XFILLER_45_484 VPWR VGND sg13g2_decap_8
X_2553_ net538 VPWR _0679_ VGND net958 net458 sg13g2_o21ai_1
X_2622_ VGND VPWR _1008_ net518 _0738_ _0737_ sg13g2_a21oi_1
X_2484_ net528 _1283_ _0622_ VPWR VGND sg13g2_nor2b_1
X_3105_ net203 VGND VPWR net762 controller.extended_cond.opcode\[0\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
X_3036_ net52 VGND VPWR net412 controller.inst_mem.mem_data\[140\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_23_123 VPWR VGND sg13g2_fill_1
XFILLER_42_498 VPWR VGND sg13g2_decap_8
XFILLER_42_421 VPWR VGND sg13g2_decap_8
XFILLER_6_399 VPWR VGND sg13g2_fill_1
XFILLER_18_451 VPWR VGND sg13g2_fill_2
XFILLER_33_465 VPWR VGND sg13g2_decap_8
X_1984_ VGND VPWR _1208_ net552 _0008_ _1318_ sg13g2_a21oi_1
X_3193__180 VPWR VGND net180 sg13g2_tiehi
X_2467_ _0608_ net457 net8 _0591_ net468 VPWR VGND sg13g2_a22oi_1
X_2536_ VGND VPWR _0662_ _0663_ _0163_ _0664_ sg13g2_a21oi_1
X_2605_ _0719_ VPWR _0721_ VGND net490 net489 sg13g2_o21ai_1
X_2398_ _0541_ net525 controller.extended_then_action\[4\] net512 controller.inst_mem.mem_data\[168\]
+ VPWR VGND sg13g2_a22oi_1
X_3011__102 VPWR VGND net102 sg13g2_tiehi
X_3019_ net86 VGND VPWR net363 controller.inst_mem.mem_data\[123\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_2
X_3029__66 VPWR VGND net66 sg13g2_tiehi
X_3092__229 VPWR VGND net229 sg13g2_tiehi
X_3061__291 VPWR VGND net291 sg13g2_tiehi
X_3172__264 VPWR VGND net264 sg13g2_tiehi
XFILLER_19_204 VPWR VGND sg13g2_fill_1
X_2321_ _0467_ net1 _0448_ VPWR VGND sg13g2_nand2b_1
XFILLER_6_163 VPWR VGND sg13g2_fill_1
X_2183_ net638 VPWR _0367_ VGND controller.inst_mem.mem_data\[189\] net573 sg13g2_o21ai_1
X_2252_ VGND VPWR _1074_ net598 _0142_ _0401_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_25 VPWR VGND uio_oe[2] sg13g2_tielo
X_1967_ net643 VPWR _1310_ VGND controller.inst_mem.mem_data\[81\] net586 sg13g2_o21ai_1
X_1898_ VPWR _1249_ _1248_ VGND sg13g2_inv_1
X_2519_ VPWR VGND net954 net462 net482 controller.alu_buffer.buffer\[11\] _0650_ net471
+ sg13g2_a221oi_1
Xheichips25_can_lehmann_fsm_36 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_16_207 VPWR VGND sg13g2_fill_2
XFILLER_12_479 VPWR VGND sg13g2_fill_2
Xhold6 _0064_ VPWR VGND net333 sg13g2_dlygate4sd3_1
XFILLER_47_387 VPWR VGND sg13g2_decap_8
X_2870_ VGND VPWR _1034_ net612 _0235_ _0926_ sg13g2_a21oi_1
X_1683_ VPWR _1034_ net818 VGND sg13g2_inv_1
Xclkbuf_leaf_10_clk clknet_3_3__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
Xhold417 _0158_ VPWR VGND net964 sg13g2_dlygate4sd3_1
X_1752_ VPWR _1103_ net682 VGND sg13g2_inv_1
Xhold406 _0167_ VPWR VGND net953 sg13g2_dlygate4sd3_1
XFILLER_7_450 VPWR VGND sg13g2_fill_2
X_1821_ VPWR _1172_ net746 VGND sg13g2_inv_1
X_3186__208 VPWR VGND net208 sg13g2_tiehi
Xhold428 controller.alu_buffer.buffer\[11\] VPWR VGND net975 sg13g2_dlygate4sd3_1
Xhold439 controller.inst_mem.addr\[2\] VPWR VGND net986 sg13g2_dlygate4sd3_1
X_2304_ VPWR VGND controller.inst_mem.mem_data\[67\] _0449_ net506 controller.inst_mem.mem_data\[163\]
+ _0450_ net510 sg13g2_a221oi_1
X_2235_ net656 VPWR _0393_ VGND controller.extended_then_action\[3\] net608 sg13g2_o21ai_1
X_2097_ net660 VPWR _0324_ VGND controller.inst_mem.mem_data\[146\] net615 sg13g2_o21ai_1
X_2166_ VGND VPWR _1117_ net559 _0099_ _0358_ sg13g2_a21oi_1
X_2999_ net126 VGND VPWR net866 controller.inst_mem.mem_data\[103\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_12_254 VPWR VGND sg13g2_fill_1
X_2020_ VGND VPWR _1190_ net581 _0026_ _1336_ sg13g2_a21oi_1
X_2853_ net658 VPWR _0918_ VGND net344 net612 sg13g2_o21ai_1
X_2922_ VGND VPWR _1008_ net591 _0261_ _0952_ sg13g2_a21oi_1
X_2784_ VGND VPWR net818 net453 _0874_ _0873_ sg13g2_a21oi_1
Xhold203 controller.inst_mem.mem_data\[46\] VPWR VGND net750 sg13g2_dlygate4sd3_1
X_1735_ VPWR _1086_ net943 VGND sg13g2_inv_1
X_1666_ VPWR _1017_ net853 VGND sg13g2_inv_1
Xhold258 controller.inst_mem.mem_data\[105\] VPWR VGND net805 sg13g2_dlygate4sd3_1
Xhold225 _0072_ VPWR VGND net772 sg13g2_dlygate4sd3_1
Xhold247 controller.inst_mem.mem_data\[158\] VPWR VGND net794 sg13g2_dlygate4sd3_1
Xhold236 controller.inst_mem.extended_word\[23\] VPWR VGND net783 sg13g2_dlygate4sd3_1
Xhold214 controller.inst_mem.extended_word\[8\] VPWR VGND net761 sg13g2_dlygate4sd3_1
X_1804_ VPWR _1155_ net330 VGND sg13g2_inv_1
Xhold269 controller.inst_mem.mem_data\[99\] VPWR VGND net816 sg13g2_dlygate4sd3_1
X_3198_ net151 VGND VPWR net373 controller.const_data\[13\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2218_ VGND VPWR _1091_ net557 _0125_ _0384_ sg13g2_a21oi_1
X_2149_ net653 VPWR _0350_ VGND controller.inst_mem.mem_data\[172\] net601 sg13g2_o21ai_1
XFILLER_49_438 VPWR VGND sg13g2_decap_8
X_3121_ net171 VGND VPWR net377 controller.extended_state\[1\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_3052_ net309 VGND VPWR net704 controller.inst_mem.mem_data\[156\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_2003_ net651 VPWR _1328_ VGND controller.inst_mem.mem_data\[99\] net601 sg13g2_o21ai_1
X_2836_ VGND VPWR _1051_ net571 _0218_ _0909_ sg13g2_a21oi_1
X_2905_ net638 VPWR _0944_ VGND net664 net574 sg13g2_o21ai_1
X_2698_ net541 VPWR _0806_ VGND net896 net444 sg13g2_o21ai_1
X_2767_ VGND VPWR _1273_ _0859_ _0860_ net452 sg13g2_a21oi_1
X_1649_ VPWR _1000_ net807 VGND sg13g2_inv_1
X_1718_ VPWR _1069_ net533 VGND sg13g2_inv_1
Xfanout524 net526 net524 VPWR VGND sg13g2_buf_8
Xfanout513 _1217_ net513 VPWR VGND sg13g2_buf_8
Xfanout502 net505 net502 VPWR VGND sg13g2_buf_8
X_3168__280 VPWR VGND net280 sg13g2_tiehi
Xfanout579 net580 net579 VPWR VGND sg13g2_buf_8
Xfanout557 net558 net557 VPWR VGND sg13g2_buf_8
Xfanout546 net547 net546 VPWR VGND sg13g2_buf_8
Xfanout535 net536 net535 VPWR VGND sg13g2_buf_8
Xfanout568 net624 net568 VPWR VGND sg13g2_buf_8
XFILLER_26_154 VPWR VGND sg13g2_fill_1
X_3071__271 VPWR VGND net271 sg13g2_tiehi
XFILLER_45_463 VPWR VGND sg13g2_decap_8
X_2483_ VPWR VGND net980 net463 net483 net977 _0621_ net472 sg13g2_a221oi_1
X_2552_ _0678_ _0677_ net466 net455 controller.alu_buffer.buffer\[9\] VPWR VGND sg13g2_a22oi_1
X_2621_ VGND VPWR controller.inst_mem.mem_data\[196\] net504 _0737_ _0736_ sg13g2_a21oi_1
X_3104_ net205 VGND VPWR _0127_ controller.inst_mem.extended_word\[8\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_3035_ net54 VGND VPWR net356 controller.inst_mem.mem_data\[139\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
XFILLER_36_496 VPWR VGND sg13g2_decap_8
X_2983__158 VPWR VGND net158 sg13g2_tiehi
X_3124__161 VPWR VGND net161 sg13g2_tiehi
X_2819_ net636 VPWR _0901_ VGND controller.const_data\[2\] net570 sg13g2_o21ai_1
XFILLER_3_507 VPWR VGND sg13g2_fill_1
XFILLER_42_477 VPWR VGND sg13g2_decap_8
XFILLER_10_352 VPWR VGND sg13g2_fill_1
XFILLER_20_105 VPWR VGND sg13g2_fill_2
X_2604_ controller.extended_then_action\[1\] net490 net489 _0720_ VPWR VGND sg13g2_or3_1
X_1983_ net629 VPWR _1318_ VGND controller.inst_mem.mem_data\[89\] net552 sg13g2_o21ai_1
XFILLER_20_116 VPWR VGND sg13g2_fill_1
X_2466_ VGND VPWR _0561_ _0607_ _0581_ net485 sg13g2_a21oi_2
X_2535_ net538 VPWR _0664_ VGND net950 net459 sg13g2_o21ai_1
X_3018_ net88 VGND VPWR _0041_ controller.inst_mem.mem_data\[122\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_1
X_2397_ VPWR VGND controller.inst_mem.mem_data\[144\] net518 net520 controller.inst_mem.mem_data\[72\]
+ _0540_ net507 sg13g2_a221oi_1
X_3138__105 VPWR VGND net105 sg13g2_tiehi
X_2320_ _0466_ _0463_ _0464_ VPWR VGND sg13g2_nand2_1
XFILLER_2_392 VPWR VGND sg13g2_fill_2
XFILLER_2_381 VPWR VGND sg13g2_fill_1
X_2251_ net648 VPWR _0401_ VGND controller.inst_mem.extended_word\[23\] net593 sg13g2_o21ai_1
X_2182_ VGND VPWR _1109_ net565 _0107_ _0366_ sg13g2_a21oi_1
X_1966_ net6 net5 _1309_ VPWR VGND sg13g2_and2_1
Xheichips25_can_lehmann_fsm_26 VPWR VGND uio_oe[3] sg13g2_tielo
Xheichips25_can_lehmann_fsm_37 VPWR VGND uio_out[6] sg13g2_tielo
X_1897_ VGND VPWR _1023_ net514 _1248_ _1247_ sg13g2_a21oi_1
X_2449_ net529 controller.alu_buffer.buffer\[3\] _0592_ VPWR VGND sg13g2_xor2_1
X_2518_ VGND VPWR _0646_ _0648_ _0160_ _0649_ sg13g2_a21oi_1
XFILLER_44_506 VPWR VGND sg13g2_fill_2
XFILLER_47_366 VPWR VGND sg13g2_decap_8
XFILLER_47_344 VPWR VGND sg13g2_fill_1
Xhold7 controller.inst_mem.extended_word\[4\] VPWR VGND net334 sg13g2_dlygate4sd3_1
X_1820_ VPWR _1171_ net382 VGND sg13g2_inv_1
X_1682_ VPWR _1033_ net396 VGND sg13g2_inv_1
Xhold429 _0160_ VPWR VGND net976 sg13g2_dlygate4sd3_1
X_3016__92 VPWR VGND net92 sg13g2_tiehi
Xhold407 controller.alu_buffer.buffer\[13\] VPWR VGND net954 sg13g2_dlygate4sd3_1
X_1751_ VPWR _1102_ net400 VGND sg13g2_inv_1
X_3031__62 VPWR VGND net62 sg13g2_tiehi
Xhold418 controller.alu_buffer.buffer\[16\] VPWR VGND net965 sg13g2_dlygate4sd3_1
X_3231__170 VPWR VGND net170 sg13g2_tiehi
X_2234_ VGND VPWR _1083_ net607 _0133_ _0392_ sg13g2_a21oi_1
X_2303_ controller.extended_cond.opcode\[2\] net523 _0449_ VPWR VGND sg13g2_and2_1
X_2165_ net630 VPWR _0358_ VGND net398 net559 sg13g2_o21ai_1
XFILLER_17_0 VPWR VGND sg13g2_fill_2
X_2096_ VGND VPWR _1152_ net615 _0064_ _0323_ sg13g2_a21oi_1
X_1949_ controller.alu_buffer.buffer\[11\] _1290_ _1293_ _1296_ VGND VPWR _1295_ sg13g2_nor4_2
X_2998_ net128 VGND VPWR net861 controller.inst_mem.mem_data\[102\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
XFILLER_29_300 VPWR VGND sg13g2_fill_2
X_3238__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_4_432 VPWR VGND sg13g2_fill_2
XFILLER_47_196 VPWR VGND sg13g2_fill_1
X_2852_ VGND VPWR _1043_ net578 _0226_ _0917_ sg13g2_a21oi_1
X_2783_ VGND VPWR _1275_ _0872_ _0873_ net453 sg13g2_a21oi_1
X_3081__251 VPWR VGND net251 sg13g2_tiehi
X_1803_ VPWR _1154_ net368 VGND sg13g2_inv_1
X_2921_ net646 VPWR _0952_ VGND controller.inst_mem.mem_data\[53\] net591 sg13g2_o21ai_1
X_1734_ VPWR _1085_ net885 VGND sg13g2_inv_1
X_1665_ VPWR _1016_ net693 VGND sg13g2_inv_1
Xhold237 controller.inst_mem.mem_data\[86\] VPWR VGND net784 sg13g2_dlygate4sd3_1
Xhold226 controller.inst_mem.mem_data\[128\] VPWR VGND net773 sg13g2_dlygate4sd3_1
Xhold248 _0078_ VPWR VGND net795 sg13g2_dlygate4sd3_1
Xhold204 controller.extended_state\[1\] VPWR VGND net751 sg13g2_dlygate4sd3_1
Xhold215 _0128_ VPWR VGND net762 sg13g2_dlygate4sd3_1
Xhold259 controller.inst_mem.mem_data\[146\] VPWR VGND net806 sg13g2_dlygate4sd3_1
X_3197_ net159 VGND VPWR _0220_ controller.const_data\[12\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2217_ net628 VPWR _0384_ VGND net701 net557 sg13g2_o21ai_1
XFILLER_26_358 VPWR VGND sg13g2_fill_1
X_3008__108 VPWR VGND net108 sg13g2_tiehi
X_2079_ net629 VPWR _0315_ VGND net351 net558 sg13g2_o21ai_1
X_2148_ VGND VPWR _1126_ net603 _0090_ _0349_ sg13g2_a21oi_1
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_39_54 VPWR VGND sg13g2_fill_2
X_2993__138 VPWR VGND net138 sg13g2_tiehi
X_3058__297 VPWR VGND net297 sg13g2_tiehi
XFILLER_44_111 VPWR VGND sg13g2_fill_1
XFILLER_39_76 VPWR VGND sg13g2_fill_2
XFILLER_17_303 VPWR VGND sg13g2_fill_1
X_3147__69 VPWR VGND net69 sg13g2_tiehi
X_3051_ net311 VGND VPWR _0074_ controller.inst_mem.mem_data\[155\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_3120_ net173 VGND VPWR _0143_ controller.extended_state\[0\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
X_2002_ VGND VPWR _1199_ net619 _0017_ _1327_ sg13g2_a21oi_1
X_2835_ net636 VPWR _0909_ VGND controller.const_data\[10\] net571 sg13g2_o21ai_1
X_2766_ _0859_ net932 _1272_ VPWR VGND sg13g2_nand2_1
X_2904_ VGND VPWR _1017_ net575 _0252_ _0943_ sg13g2_a21oi_1
X_2697_ _0805_ net448 _0804_ _0767_ net788 VPWR VGND sg13g2_a22oi_1
X_1648_ VPWR _0999_ net864 VGND sg13g2_inv_1
Xfanout514 net516 net514 VPWR VGND sg13g2_buf_8
Xfanout536 net985 net536 VPWR VGND sg13g2_buf_8
X_1717_ _1068_ net531 VPWR VGND sg13g2_inv_2
Xfanout547 net554 net547 VPWR VGND sg13g2_buf_8
Xfanout503 net505 net503 VPWR VGND sg13g2_buf_8
Xfanout525 net526 net525 VPWR VGND sg13g2_buf_8
Xfanout569 net570 net569 VPWR VGND sg13g2_buf_8
XFILLER_39_494 VPWR VGND sg13g2_decap_8
X_3249_ net163 VGND VPWR _0272_ controller.inst_mem.mem_data\[64\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
Xfanout558 net568 net558 VPWR VGND sg13g2_buf_8
XFILLER_22_372 VPWR VGND sg13g2_fill_2
X_3175__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_45_442 VPWR VGND sg13g2_decap_8
XFILLER_17_155 VPWR VGND sg13g2_fill_2
X_2620_ _0734_ _0735_ _0733_ _0736_ VPWR VGND sg13g2_nand3_1
X_2482_ VGND VPWR _0618_ _0619_ _0153_ _0620_ sg13g2_a21oi_1
X_2551_ _0669_ net958 _0677_ VPWR VGND sg13g2_xor2_1
X_3103_ net207 VGND VPWR net702 controller.inst_mem.extended_word\[7\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_3034_ net56 VGND VPWR net352 controller.inst_mem.mem_data\[138\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
XFILLER_36_475 VPWR VGND sg13g2_decap_8
X_2818_ VGND VPWR _1060_ net570 _0209_ _0900_ sg13g2_a21oi_1
X_2749_ net543 VPWR _0846_ VGND net890 net477 sg13g2_o21ai_1
X_3131__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_42_456 VPWR VGND sg13g2_decap_8
X_3140__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_45_250 VPWR VGND sg13g2_fill_1
XFILLER_33_434 VPWR VGND sg13g2_fill_1
X_1982_ VGND VPWR _1209_ net546 _0007_ _1317_ sg13g2_a21oi_1
X_2534_ _0663_ net455 net527 net471 controller.alu_buffer.buffer\[13\] VPWR VGND sg13g2_a22oi_1
X_2603_ _0718_ VPWR _0719_ VGND controller.inst_mem.mem_data\[51\] net491 sg13g2_o21ai_1
XFILLER_47_0 VPWR VGND sg13g2_fill_2
X_2465_ _0605_ _0606_ _0150_ VPWR VGND sg13g2_nor2_1
X_2396_ _0539_ net495 controller.inst_mem.mem_data\[96\] net503 controller.inst_mem.mem_data\[192\]
+ VPWR VGND sg13g2_a22oi_1
X_3017_ net90 VGND VPWR _0040_ controller.inst_mem.mem_data\[121\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_1
XFILLER_22_35 VPWR VGND sg13g2_fill_1
XFILLER_42_286 VPWR VGND sg13g2_fill_2
XFILLER_15_412 VPWR VGND sg13g2_fill_1
X_3257__190 VPWR VGND net190 sg13g2_tiehi
X_2250_ VGND VPWR _1075_ net598 _0141_ _0400_ sg13g2_a21oi_1
X_2181_ net638 VPWR _0366_ VGND net438 net572 sg13g2_o21ai_1
X_1965_ net22 _1307_ _1308_ VPWR VGND sg13g2_nand2_1
Xheichips25_can_lehmann_fsm_27 VPWR VGND uio_oe[4] sg13g2_tielo
X_2517_ net538 VPWR _0649_ VGND net975 net459 sg13g2_o21ai_1
X_3091__231 VPWR VGND net231 sg13g2_tiehi
X_1896_ VGND VPWR controller.inst_mem.mem_data\[61\] net506 _1247_ _1246_ sg13g2_a21oi_1
Xheichips25_can_lehmann_fsm_38 VPWR VGND uio_out[7] sg13g2_tielo
X_2448_ _0591_ net530 net971 VPWR VGND sg13g2_xnor2_1
X_2379_ _0522_ VPWR _0523_ VGND net800 net491 sg13g2_o21ai_1
XFILLER_33_89 VPWR VGND sg13g2_fill_1
XFILLER_3_168 VPWR VGND sg13g2_fill_2
XFILLER_35_507 VPWR VGND sg13g2_fill_1
Xhold8 _0124_ VPWR VGND net335 sg13g2_dlygate4sd3_1
X_3068__277 VPWR VGND net277 sg13g2_tiehi
X_1750_ VPWR _1101_ net790 VGND sg13g2_inv_1
X_1681_ VPWR _1032_ net822 VGND sg13g2_inv_1
Xhold408 _0162_ VPWR VGND net955 sg13g2_dlygate4sd3_1
Xhold419 _0165_ VPWR VGND net966 sg13g2_dlygate4sd3_1
XFILLER_38_345 VPWR VGND sg13g2_fill_2
X_2233_ net655 VPWR _0392_ VGND net685 net607 sg13g2_o21ai_1
X_2164_ VGND VPWR _1118_ net584 _0098_ _0357_ sg13g2_a21oi_1
X_2302_ _0448_ _0445_ _0447_ net515 _1018_ VPWR VGND sg13g2_a22oi_1
XFILLER_21_201 VPWR VGND sg13g2_fill_1
X_2095_ net660 VPWR _0323_ VGND controller.inst_mem.mem_data\[145\] net615 sg13g2_o21ai_1
X_1948_ controller.alu_buffer.buffer\[19\] controller.alu_buffer.buffer\[18\] controller.alu_buffer.buffer\[17\]
+ controller.alu_buffer.buffer\[16\] _1295_ VPWR VGND sg13g2_or4_1
X_1879_ net533 net536 _1230_ VPWR VGND sg13g2_nor2_1
X_2997_ net130 VGND VPWR net837 controller.inst_mem.mem_data\[101\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_0_105 VPWR VGND sg13g2_fill_1
XFILLER_12_212 VPWR VGND sg13g2_fill_2
X_2920_ VGND VPWR _1009_ net588 _0260_ _0951_ sg13g2_a21oi_1
X_2851_ net640 VPWR _0917_ VGND net409 net576 sg13g2_o21ai_1
X_2782_ _0872_ net907 _1274_ VPWR VGND sg13g2_nand2b_1
X_1733_ VPWR _1084_ net858 VGND sg13g2_inv_1
X_1802_ VPWR _1153_ net781 VGND sg13g2_inv_1
Xhold227 controller.const_data\[5\] VPWR VGND net774 sg13g2_dlygate4sd3_1
X_1664_ VPWR _1015_ net664 VGND sg13g2_inv_1
Xhold238 _0006_ VPWR VGND net785 sg13g2_dlygate4sd3_1
Xhold249 controller.inst_mem.mem_data\[85\] VPWR VGND net796 sg13g2_dlygate4sd3_1
Xhold216 controller.inst_mem.mem_data\[114\] VPWR VGND net763 sg13g2_dlygate4sd3_1
Xhold205 _0145_ VPWR VGND net752 sg13g2_dlygate4sd3_1
X_3196_ net167 VGND VPWR _0219_ controller.const_data\[11\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2216_ VGND VPWR _1092_ net561 _0124_ _0383_ sg13g2_a21oi_1
X_3265_ net270 VGND VPWR _0288_ controller.inst_mem.mem_data\[80\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_2147_ net651 VPWR _0349_ VGND net744 net603 sg13g2_o21ai_1
X_2078_ VGND VPWR _1161_ net552 _0055_ _0314_ sg13g2_a21oi_1
XFILLER_32_318 VPWR VGND sg13g2_fill_1
X_3256__222 VPWR VGND net222 sg13g2_tiehi
XFILLER_48_484 VPWR VGND sg13g2_decap_8
X_3050_ net313 VGND VPWR _0073_ controller.inst_mem.mem_data\[154\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_2001_ net661 VPWR _1327_ VGND controller.inst_mem.mem_data\[98\] net619 sg13g2_o21ai_1
X_2903_ net639 VPWR _0943_ VGND net693 net575 sg13g2_o21ai_1
XFILLER_23_318 VPWR VGND sg13g2_fill_2
X_2834_ VGND VPWR _1052_ net571 _0217_ _0908_ sg13g2_a21oi_1
X_2765_ VGND VPWR net477 _0857_ _0198_ _0858_ sg13g2_a21oi_1
X_2696_ _0804_ net896 _0411_ VPWR VGND sg13g2_xnor2_1
X_1716_ VPWR _1067_ net971 VGND sg13g2_inv_1
Xfanout537 net542 net537 VPWR VGND sg13g2_buf_8
Xfanout559 net561 net559 VPWR VGND sg13g2_buf_8
X_1647_ VPWR _0998_ net758 VGND sg13g2_inv_1
Xfanout548 net549 net548 VPWR VGND sg13g2_buf_8
Xfanout526 _1229_ net526 VPWR VGND sg13g2_buf_8
Xfanout504 net505 net504 VPWR VGND sg13g2_buf_8
Xfanout515 net516 net515 VPWR VGND sg13g2_buf_8
XFILLER_39_473 VPWR VGND sg13g2_decap_8
X_3179_ net236 VGND VPWR net908 controller.counter2.counter_1\[10\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
X_3248_ net182 VGND VPWR net759 controller.inst_mem.mem_data\[63\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_41_45 VPWR VGND sg13g2_fill_2
XFILLER_45_421 VPWR VGND sg13g2_decap_8
XFILLER_45_498 VPWR VGND sg13g2_decap_8
XFILLER_32_126 VPWR VGND sg13g2_fill_2
X_3182__224 VPWR VGND net224 sg13g2_tiehi
X_2550_ controller.alu_buffer.buffer\[17\] controller.alu_buffer.buffer\[16\] _1294_
+ _0676_ VPWR VGND sg13g2_nor3_1
X_2481_ net539 VPWR _0620_ VGND net977 net460 sg13g2_o21ai_1
X_3050__313 VPWR VGND net313 sg13g2_tiehi
X_3161__308 VPWR VGND net308 sg13g2_tiehi
XFILLER_36_454 VPWR VGND sg13g2_decap_8
X_3102_ net209 VGND VPWR _0125_ controller.inst_mem.extended_word\[6\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_3033_ net58 VGND VPWR _0056_ controller.inst_mem.mem_data\[137\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_2817_ net636 VPWR _0900_ VGND controller.const_data\[1\] net570 sg13g2_o21ai_1
X_2679_ VPWR VGND net11 net446 _0774_ net419 _0791_ net479 sg13g2_a221oi_1
X_2748_ VGND VPWR net344 net451 _0845_ _0844_ sg13g2_a21oi_1
XFILLER_11_48 VPWR VGND sg13g2_fill_2
XFILLER_42_435 VPWR VGND sg13g2_decap_8
XFILLER_6_303 VPWR VGND sg13g2_fill_2
XFILLER_33_479 VPWR VGND sg13g2_decap_8
X_3258__147 VPWR VGND net147 sg13g2_tiehi
X_2982__160 VPWR VGND net160 sg13g2_tiehi
X_1981_ net626 VPWR _1317_ VGND net370 net551 sg13g2_o21ai_1
X_2533_ VPWR VGND net466 net461 _0661_ net922 _0662_ net482 sg13g2_a221oi_1
X_3078__257 VPWR VGND net257 sg13g2_tiehi
X_2602_ _0715_ _0716_ _0714_ _0718_ VPWR VGND _0717_ sg13g2_nand4_1
X_2464_ net539 VPWR _0606_ VGND net971 _0596_ sg13g2_o21ai_1
X_2395_ _0538_ controller.inst_mem.mem_data\[120\] net499 VPWR VGND sg13g2_nand2_1
X_3016_ net92 VGND VPWR _0039_ controller.inst_mem.mem_data\[120\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_31_clk clknet_3_4__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
XFILLER_30_438 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_22_clk clknet_3_7__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
X_2180_ VGND VPWR _1110_ net564 _0106_ _0365_ sg13g2_a21oi_1
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_1964_ _1308_ _1258_ controller.alu_buffer.buffer\[7\] _1257_ net532 VPWR VGND sg13g2_a22oi_1
X_1895_ _1244_ _1245_ _1243_ _1246_ VPWR VGND sg13g2_nand3_1
X_2447_ _0590_ _0588_ _0589_ VPWR VGND sg13g2_xnor2_1
X_2516_ _0648_ _0647_ net467 net456 controller.alu_buffer.buffer\[3\] VPWR VGND sg13g2_a22oi_1
Xheichips25_can_lehmann_fsm_28 VPWR VGND uio_oe[5] sg13g2_tielo
X_2378_ _0519_ _0520_ _0518_ _0522_ VPWR VGND _0521_ sg13g2_nand4_1
Xhold9 controller.inst_mem.mem_data\[168\] VPWR VGND net336 sg13g2_dlygate4sd3_1
X_1680_ VPWR _1031_ net440 VGND sg13g2_inv_1
Xhold409 controller.alu_buffer.buffer\[22\] VPWR VGND net956 sg13g2_dlygate4sd3_1
XFILLER_7_497 VPWR VGND sg13g2_fill_1
X_2301_ net515 _0441_ _0444_ _0446_ _0447_ VPWR VGND sg13g2_nor4_1
X_2232_ VGND VPWR _1084_ net572 _0132_ _0391_ sg13g2_a21oi_1
X_2163_ net642 VPWR _0357_ VGND net706 net581 sg13g2_o21ai_1
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2094_ VGND VPWR _1153_ net608 _0063_ _0322_ sg13g2_a21oi_1
XFILLER_0_72 VPWR VGND sg13g2_fill_1
X_1947_ VGND VPWR _1294_ _1293_ _1291_ sg13g2_or2_1
X_1878_ _1229_ net532 net533 net536 VPWR VGND sg13g2_and3_1
X_2996_ net132 VGND VPWR net817 controller.inst_mem.mem_data\[100\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
XFILLER_44_338 VPWR VGND sg13g2_fill_2
X_3178__240 VPWR VGND net240 sg13g2_tiehi
X_2850_ VGND VPWR _1044_ net576 _0225_ _0916_ sg13g2_a21oi_1
XFILLER_31_500 VPWR VGND sg13g2_decap_8
X_3157__324 VPWR VGND net324 sg13g2_tiehi
X_2781_ VGND VPWR net478 _0870_ _0201_ _0871_ sg13g2_a21oi_1
X_1663_ VPWR _1014_ net750 VGND sg13g2_inv_1
X_1732_ VPWR _1083_ net728 VGND sg13g2_inv_1
Xhold206 controller.inst_mem.mem_data\[169\] VPWR VGND net753 sg13g2_dlygate4sd3_1
Xhold217 _0034_ VPWR VGND net764 sg13g2_dlygate4sd3_1
X_1801_ VPWR _1152_ net332 VGND sg13g2_inv_1
Xhold228 controller.inst_mem.mem_data\[107\] VPWR VGND net775 sg13g2_dlygate4sd3_1
X_3264_ net206 VGND VPWR _0287_ controller.inst_mem.mem_data\[79\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_2
Xhold239 controller.inst_mem.mem_data\[52\] VPWR VGND net786 sg13g2_dlygate4sd3_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
X_3195_ net172 VGND VPWR net391 controller.const_data\[10\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_26_305 VPWR VGND sg13g2_fill_2
X_2146_ VGND VPWR _1127_ net619 _0089_ _0348_ sg13g2_a21oi_1
X_2215_ net630 VPWR _0383_ VGND controller.inst_mem.extended_word\[5\] net556 sg13g2_o21ai_1
X_2077_ net629 VPWR _0314_ VGND net435 net552 sg13g2_o21ai_1
X_3197__159 VPWR VGND net159 sg13g2_tiehi
X_2979_ net166 VGND VPWR net678 controller.inst_mem.mem_data\[83\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_3134__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_44_179 VPWR VGND sg13g2_fill_2
X_3106__201 VPWR VGND net201 sg13g2_tiehi
XFILLER_48_463 VPWR VGND sg13g2_decap_8
X_2000_ VGND VPWR _1200_ net618 _0016_ _1326_ sg13g2_a21oi_1
X_2833_ net637 VPWR _0908_ VGND net390 net571 sg13g2_o21ai_1
X_3007__110 VPWR VGND net110 sg13g2_tiehi
X_2902_ VGND VPWR _1018_ net563 _0251_ _0942_ sg13g2_a21oi_1
X_2764_ net543 VPWR _0858_ VGND net888 net477 sg13g2_o21ai_1
X_1715_ VPWR _1066_ controller.alu_buffer.buffer\[5\] VGND sg13g2_inv_1
X_2695_ VPWR VGND _0803_ _0503_ _0802_ _1063_ _0183_ net447 sg13g2_a221oi_1
X_2992__140 VPWR VGND net140 sg13g2_tiehi
X_1646_ VPWR _0997_ net862 VGND sg13g2_inv_1
XFILLER_39_452 VPWR VGND sg13g2_decap_8
Xfanout527 net982 net527 VPWR VGND sg13g2_buf_8
Xfanout538 net542 net538 VPWR VGND sg13g2_buf_8
X_3088__237 VPWR VGND net237 sg13g2_tiehi
X_3247_ net198 VGND VPWR _0270_ controller.inst_mem.mem_data\[62\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
Xfanout549 net550 net549 VPWR VGND sg13g2_buf_8
Xfanout505 _1222_ net505 VPWR VGND sg13g2_buf_8
Xfanout516 _1231_ net516 VPWR VGND sg13g2_buf_8
X_3178_ net240 VGND VPWR net902 controller.counter2.counter_1\[9\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
X_2129_ net632 VPWR _0340_ VGND controller.inst_mem.mem_data\[162\] net562 sg13g2_o21ai_1
XFILLER_45_400 VPWR VGND sg13g2_decap_8
XFILLER_45_477 VPWR VGND sg13g2_decap_8
XFILLER_17_179 VPWR VGND sg13g2_fill_1
X_2480_ _0619_ net457 net10 net472 net529 VPWR VGND sg13g2_a22oi_1
X_3101_ net211 VGND VPWR net335 controller.inst_mem.extended_word\[5\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_3143__85 VPWR VGND net85 sg13g2_tiehi
X_3032_ net60 VGND VPWR _0055_ controller.inst_mem.mem_data\[136\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_2816_ VGND VPWR _1061_ net580 _0208_ _0899_ sg13g2_a21oi_1
X_2678_ net448 VPWR _0790_ VGND _0408_ _0789_ sg13g2_o21ai_1
X_2747_ VGND VPWR _1270_ _0843_ _0844_ net451 sg13g2_a21oi_1
X_1629_ VPWR _0980_ net414 VGND sg13g2_inv_1
XFILLER_14_116 VPWR VGND sg13g2_fill_1
XFILLER_22_171 VPWR VGND sg13g2_fill_2
X_1980_ VGND VPWR _1210_ net548 _0006_ _1316_ sg13g2_a21oi_1
X_3038__48 VPWR VGND net48 sg13g2_tiehi
X_2463_ VPWR VGND net530 _0604_ net484 _1067_ _0605_ net468 sg13g2_a221oi_1
X_2532_ _0656_ net950 _0661_ VPWR VGND sg13g2_xor2_1
X_2601_ _0717_ net500 controller.inst_mem.mem_data\[123\] net504 controller.inst_mem.mem_data\[195\]
+ VPWR VGND sg13g2_a22oi_1
X_3015_ net94 VGND VPWR net769 controller.inst_mem.mem_data\[119\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_2394_ _0528_ _0536_ net486 _0537_ VPWR VGND sg13g2_nand3_1
XFILLER_47_506 VPWR VGND sg13g2_fill_2
XFILLER_27_241 VPWR VGND sg13g2_fill_1
X_3220__258 VPWR VGND net258 sg13g2_tiehi
X_3114__185 VPWR VGND net185 sg13g2_tiehi
X_1894_ VPWR VGND controller.inst_mem.mem_data\[133\] net514 net519 controller.inst_mem.mem_data\[109\]
+ _1245_ net498 sg13g2_a221oi_1
X_1963_ _1307_ controller.alu_buffer.buffer\[23\] _1260_ VPWR VGND sg13g2_nand2_1
X_2446_ net528 controller.alu_buffer.buffer\[5\] _0589_ VPWR VGND sg13g2_xor2_1
X_2515_ _0647_ net975 _1290_ VPWR VGND sg13g2_xnor2_1
Xheichips25_can_lehmann_fsm_29 VPWR VGND uio_oe[6] sg13g2_tielo
X_2377_ VGND VPWR controller.inst_mem.mem_data\[154\] net511 _0521_ net517 sg13g2_a21oi_1
X_2231_ net638 VPWR _0391_ VGND net728 net572 sg13g2_o21ai_1
X_2300_ _0442_ VPWR _0446_ VGND _1134_ _1218_ sg13g2_o21ai_1
X_2162_ VGND VPWR _1119_ net585 _0097_ _0356_ sg13g2_a21oi_1
X_3047__319 VPWR VGND net319 sg13g2_tiehi
X_2093_ net660 VPWR _0322_ VGND net332 net616 sg13g2_o21ai_1
X_2995_ net134 VGND VPWR net709 controller.inst_mem.mem_data\[99\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_1946_ _1293_ _1064_ _1292_ VPWR VGND sg13g2_nand2_1
X_1877_ _1228_ net494 controller.inst_mem.mem_data\[87\] net498 controller.inst_mem.mem_data\[111\]
+ VPWR VGND sg13g2_a22oi_1
X_2429_ _0571_ VPWR _0572_ VGND net490 net489 sg13g2_o21ai_1
X_3098__217 VPWR VGND net217 sg13g2_tiehi
X_3013__98 VPWR VGND net98 sg13g2_tiehi
X_3185__212 VPWR VGND net212 sg13g2_tiehi
X_1800_ VPWR _1151_ net679 VGND sg13g2_inv_1
X_2780_ net543 VPWR _0871_ VGND net901 net478 sg13g2_o21ai_1
X_1662_ VPWR _1013_ net413 VGND sg13g2_inv_1
Xhold207 _0089_ VPWR VGND net754 sg13g2_dlygate4sd3_1
Xhold229 _0027_ VPWR VGND net776 sg13g2_dlygate4sd3_1
X_2979__166 VPWR VGND net166 sg13g2_tiehi
Xhold218 controller.inst_mem.mem_data\[58\] VPWR VGND net765 sg13g2_dlygate4sd3_1
X_1731_ VPWR _1082_ net685 VGND sg13g2_inv_1
X_3194_ net176 VGND VPWR _0217_ controller.const_data\[9\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2214_ VGND VPWR _1093_ net561 _0123_ _0382_ sg13g2_a21oi_1
X_3263_ net45 VGND VPWR net827 controller.inst_mem.mem_data\[78\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_2145_ net661 VPWR _0348_ VGND controller.inst_mem.mem_data\[170\] net619 sg13g2_o21ai_1
X_2076_ VGND VPWR _1162_ net550 _0054_ _0313_ sg13g2_a21oi_1
XFILLER_15_0 VPWR VGND sg13g2_fill_2
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
X_1929_ _1277_ _1274_ _1276_ VPWR VGND sg13g2_nand2_2
X_2978_ net168 VGND VPWR _0001_ controller.inst_mem.mem_data\[82\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
X_3156__39 VPWR VGND net39 sg13g2_tiehi
XFILLER_17_317 VPWR VGND sg13g2_fill_1
XFILLER_48_442 VPWR VGND sg13g2_decap_8
Xhold90 _0026_ VPWR VGND net417 sg13g2_dlygate4sd3_1
X_2832_ VGND VPWR _1053_ net570 _0216_ _0907_ sg13g2_a21oi_1
X_2763_ VGND VPWR net840 net453 _0857_ _0856_ sg13g2_a21oi_1
X_2901_ net634 VPWR _0942_ VGND controller.inst_mem.mem_data\[43\] net563 sg13g2_o21ai_1
X_2694_ VPWR VGND net14 net446 _0774_ net824 _0803_ net479 sg13g2_a221oi_1
X_1645_ VPWR _0996_ net328 VGND sg13g2_inv_1
X_1714_ VPWR _1065_ net963 VGND sg13g2_inv_1
Xfanout506 net509 net506 VPWR VGND sg13g2_buf_8
Xfanout539 net541 net539 VPWR VGND sg13g2_buf_8
Xfanout528 net961 net528 VPWR VGND sg13g2_buf_8
X_3177_ net244 VGND VPWR _0200_ controller.counter2.counter_1\[8\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_2
X_3246_ net214 VGND VPWR net808 controller.inst_mem.mem_data\[61\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
Xfanout517 net518 net517 VPWR VGND sg13g2_buf_8
XFILLER_26_147 VPWR VGND sg13g2_fill_2
X_2059_ net650 VPWR _0305_ VGND controller.inst_mem.mem_data\[127\] net596 sg13g2_o21ai_1
X_2128_ VGND VPWR _1136_ net551 _0080_ _0339_ sg13g2_a21oi_1
X_3152__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_45_456 VPWR VGND sg13g2_decap_8
X_3223__234 VPWR VGND net234 sg13g2_tiehi
X_3031_ net62 VGND VPWR net429 controller.inst_mem.mem_data\[135\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_3100_ net213 VGND VPWR _0123_ controller.inst_mem.extended_word\[4\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_36_489 VPWR VGND sg13g2_decap_8
XFILLER_23_128 VPWR VGND sg13g2_fill_1
X_2746_ _0843_ net890 _1269_ VPWR VGND sg13g2_nand2b_1
X_2815_ net637 VPWR _0899_ VGND net671 net580 sg13g2_o21ai_1
X_2677_ net944 _0407_ _0789_ VPWR VGND sg13g2_and2_1
XFILLER_39_272 VPWR VGND sg13g2_fill_1
X_3229_ net186 VGND VPWR _0252_ controller.inst_mem.mem_data\[44\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
XFILLER_10_367 VPWR VGND sg13g2_fill_2
Xhold390 _0129_ VPWR VGND net937 sg13g2_dlygate4sd3_1
XFILLER_41_481 VPWR VGND sg13g2_decap_8
X_2600_ _0716_ net496 controller.inst_mem.mem_data\[99\] net508 controller.inst_mem.mem_data\[75\]
+ VPWR VGND sg13g2_a22oi_1
X_3210__49 VPWR VGND net49 sg13g2_tiehi
X_2462_ _0604_ net460 _1061_ _0583_ _0562_ VPWR VGND sg13g2_a22oi_1
X_2531_ _1291_ _1292_ _0660_ VPWR VGND sg13g2_nor2b_1
X_2393_ _0535_ VPWR _0536_ VGND net490 net489 sg13g2_o21ai_1
X_3014_ net96 VGND VPWR _0037_ controller.inst_mem.mem_data\[118\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
XFILLER_32_481 VPWR VGND sg13g2_decap_8
X_2729_ _0828_ _0829_ _0191_ VPWR VGND sg13g2_nor2_1
XFILLER_15_404 VPWR VGND sg13g2_fill_2
XFILLER_6_179 VPWR VGND sg13g2_fill_2
XFILLER_10_197 VPWR VGND sg13g2_fill_1
XFILLER_38_507 VPWR VGND sg13g2_fill_1
X_1962_ net21 _1305_ _1306_ VPWR VGND sg13g2_nand2_2
X_1893_ _1244_ net502 controller.inst_mem.mem_data\[181\] net510 controller.inst_mem.mem_data\[157\]
+ VPWR VGND sg13g2_a22oi_1
X_2445_ net527 controller.alu_buffer.buffer\[7\] _0588_ VPWR VGND sg13g2_xor2_1
X_2514_ VPWR VGND net969 net462 net482 controller.alu_buffer.buffer\[10\] _0646_ net471
+ sg13g2_a221oi_1
X_2376_ _0520_ _0479_ controller.inst_mem.mem_data\[130\] net495 controller.inst_mem.mem_data\[82\]
+ VPWR VGND sg13g2_a22oi_1
X_2989__146 VPWR VGND net146 sg13g2_tiehi
X_3025__74 VPWR VGND net74 sg13g2_tiehi
X_3040__44 VPWR VGND net44 sg13g2_tiehi
X_2230_ VGND VPWR _1085_ net575 _0131_ _0390_ sg13g2_a21oi_1
XFILLER_46_392 VPWR VGND sg13g2_decap_8
X_2161_ net643 VPWR _0356_ VGND controller.inst_mem.mem_data\[178\] net585 sg13g2_o21ai_1
X_2092_ VGND VPWR _1154_ net588 _0062_ _0321_ sg13g2_a21oi_1
X_1945_ controller.alu_buffer.buffer\[14\] controller.alu_buffer.buffer\[13\] controller.alu_buffer.buffer\[12\]
+ _1292_ VPWR VGND sg13g2_nor3_1
X_2994_ net136 VGND VPWR net422 controller.inst_mem.mem_data\[98\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_1876_ net531 _1221_ _1227_ VPWR VGND sg13g2_nor2_1
XFILLER_29_315 VPWR VGND sg13g2_fill_1
X_2359_ VGND VPWR _1070_ _0494_ _0146_ _0504_ sg13g2_a21oi_1
X_2428_ VPWR _0571_ _0570_ VGND sg13g2_inv_1
XFILLER_44_47 VPWR VGND sg13g2_fill_1
XFILLER_20_281 VPWR VGND sg13g2_fill_1
XFILLER_35_307 VPWR VGND sg13g2_fill_2
X_3226__210 VPWR VGND net210 sg13g2_tiehi
X_3265__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_18_70 VPWR VGND sg13g2_fill_1
X_1661_ VPWR _1012_ net407 VGND sg13g2_inv_1
X_1730_ VPWR _1081_ net882 VGND sg13g2_inv_1
Xhold219 _0267_ VPWR VGND net766 sg13g2_dlygate4sd3_1
Xhold208 controller.inst_mem.mem_data\[198\] VPWR VGND net755 sg13g2_dlygate4sd3_1
X_3193_ net180 VGND VPWR _0216_ controller.const_data\[8\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2144_ VGND VPWR _1128_ net615 _0088_ _0347_ sg13g2_a21oi_1
X_2213_ net630 VPWR _0382_ VGND net334 net561 sg13g2_o21ai_1
X_3262_ net174 VGND VPWR _0285_ controller.inst_mem.mem_data\[77\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
X_2075_ net626 VPWR _0313_ VGND controller.inst_mem.mem_data\[135\] net550 sg13g2_o21ai_1
X_1928_ net883 controller.counter2.counter_1\[10\] _1276_ VPWR VGND sg13g2_nor2_1
X_1859_ VPWR _1210_ net784 VGND sg13g2_inv_1
X_2977_ net115 VGND VPWR net415 controller.inst_mem.mem_data\[81\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_25_373 VPWR VGND sg13g2_fill_2
XFILLER_48_421 VPWR VGND sg13g2_decap_8
XFILLER_48_498 VPWR VGND sg13g2_decap_8
Xhold91 controller.const_data\[16\] VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold80 controller.inst_mem.mem_data\[48\] VPWR VGND net407 sg13g2_dlygate4sd3_1
X_2900_ VGND VPWR _1019_ net563 _0250_ _0941_ sg13g2_a21oi_1
X_2831_ net637 VPWR _0907_ VGND net788 net571 sg13g2_o21ai_1
X_2762_ VGND VPWR _1272_ _0855_ _0856_ net452 sg13g2_a21oi_1
X_1713_ _1064_ net922 VPWR VGND sg13g2_inv_2
Xfanout529 net933 net529 VPWR VGND sg13g2_buf_8
X_2693_ _0802_ net449 _0801_ VPWR VGND sg13g2_nand2_1
X_1644_ VPWR _0995_ net374 VGND sg13g2_inv_1
Xfanout507 net509 net507 VPWR VGND sg13g2_buf_8
X_3146__73 VPWR VGND net73 sg13g2_tiehi
Xfanout518 _1231_ net518 VPWR VGND sg13g2_buf_8
XFILLER_39_487 VPWR VGND sg13g2_decap_8
X_3176_ net248 VGND VPWR _0199_ controller.counter2.counter_1\[7\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_2
X_3245_ net230 VGND VPWR _0268_ controller.inst_mem.mem_data\[60\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_2127_ net626 VPWR _0339_ VGND net338 net551 sg13g2_o21ai_1
X_2058_ VGND VPWR _1171_ net596 _0045_ _0304_ sg13g2_a21oi_1
XFILLER_45_435 VPWR VGND sg13g2_decap_8
X_3030_ net64 VGND VPWR net385 controller.inst_mem.mem_data\[134\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_36_468 VPWR VGND sg13g2_decap_8
X_2745_ VGND VPWR net475 _0841_ _0194_ _0842_ sg13g2_a21oi_1
X_2676_ VGND VPWR _0786_ _0787_ _0179_ _0788_ sg13g2_a21oi_1
X_2814_ VGND VPWR net474 _0897_ _0207_ _0898_ sg13g2_a21oi_1
X_3159_ net316 VGND VPWR net895 controller.counter2.counter_0\[6\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
X_3228_ net194 VGND VPWR net741 controller.inst_mem.mem_data\[43\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
XFILLER_42_449 VPWR VGND sg13g2_decap_8
X_2999__126 VPWR VGND net126 sg13g2_tiehi
Xclkbuf_leaf_34_clk clknet_3_1__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
Xhold380 _0205_ VPWR VGND net927 sg13g2_dlygate4sd3_1
Xhold391 controller.counter2.counter_0\[5\] VPWR VGND net938 sg13g2_dlygate4sd3_1
XFILLER_41_460 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_3_5__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
X_2530_ VGND VPWR _0655_ _0658_ _0162_ _0659_ sg13g2_a21oi_1
X_2461_ VPWR VGND _0553_ _0560_ _0546_ _0537_ _0603_ _0544_ sg13g2_a221oi_1
XFILLER_5_383 VPWR VGND sg13g2_fill_1
X_2392_ VPWR _0535_ _0534_ VGND sg13g2_inv_1
X_3013_ net98 VGND VPWR net674 controller.inst_mem.mem_data\[117\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_16_clk clknet_3_6__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_3037__50 VPWR VGND net50 sg13g2_tiehi
X_2659_ VPWR VGND net7 net447 _0774_ net671 _0775_ net479 sg13g2_a221oi_1
X_2728_ net541 VPWR _0829_ VGND net906 net445 sg13g2_o21ai_1
XFILLER_10_176 VPWR VGND sg13g2_fill_2
X_3188__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_12_83 VPWR VGND sg13g2_fill_1
XFILLER_37_91 VPWR VGND sg13g2_fill_1
XFILLER_33_268 VPWR VGND sg13g2_fill_1
XFILLER_33_235 VPWR VGND sg13g2_fill_2
X_1961_ _1306_ _1258_ net527 _1257_ net533 VPWR VGND sg13g2_a22oi_1
X_1892_ _1243_ net523 controller.inst_mem.extended_word\[5\] net494 controller.inst_mem.mem_data\[85\]
+ VPWR VGND sg13g2_a22oi_1
X_2513_ VGND VPWR _0643_ net934 _0159_ _0645_ sg13g2_a21oi_1
X_2444_ _0587_ controller.alu_buffer.buffer\[8\] _1287_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_5_clk clknet_3_3__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2375_ _0519_ net499 controller.inst_mem.mem_data\[106\] net503 controller.inst_mem.mem_data\[178\]
+ VPWR VGND sg13g2_a22oi_1
X_2160_ VGND VPWR _1120_ net592 _0096_ _0355_ sg13g2_a21oi_1
X_2091_ net646 VPWR _0321_ VGND controller.inst_mem.mem_data\[143\] net588 sg13g2_o21ai_1
X_2993_ net138 VGND VPWR _0016_ controller.inst_mem.mem_data\[97\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
X_1944_ VGND VPWR _1291_ _1290_ controller.alu_buffer.buffer\[11\] sg13g2_or2_1
X_1875_ net531 _1225_ _1226_ VPWR VGND sg13g2_nor2_1
X_2427_ _0569_ VPWR _0570_ VGND controller.inst_mem.mem_data\[53\] net491 sg13g2_o21ai_1
X_2289_ _0431_ _0434_ _0435_ VPWR VGND sg13g2_nor2_1
X_2358_ net545 VPWR _0504_ VGND _0494_ _0501_ sg13g2_o21ai_1
X_3046__321 VPWR VGND net321 sg13g2_tiehi
X_3237__75 VPWR VGND net75 sg13g2_tiehi
X_3252__67 VPWR VGND net67 sg13g2_tiehi
X_1660_ VPWR _1011_ net852 VGND sg13g2_inv_1
Xhold209 _0118_ VPWR VGND net756 sg13g2_dlygate4sd3_1
X_3192_ net184 VGND VPWR net716 controller.const_data\[7\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2143_ net660 VPWR _0347_ VGND controller.inst_mem.mem_data\[169\] net615 sg13g2_o21ai_1
X_2212_ VGND VPWR _1094_ net582 _0122_ _0381_ sg13g2_a21oi_1
X_3261_ net238 VGND VPWR net793 controller.inst_mem.mem_data\[76\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_2074_ VGND VPWR _1163_ net557 _0053_ _0312_ sg13g2_a21oi_1
X_1927_ _1275_ _1274_ net907 VPWR VGND sg13g2_nand2b_1
X_1858_ VPWR _1209_ net789 VGND sg13g2_inv_1
X_2976_ VGND VPWR _0981_ net594 _0288_ _0979_ sg13g2_a21oi_1
X_1789_ VPWR _1140_ net875 VGND sg13g2_inv_1
XFILLER_29_113 VPWR VGND sg13g2_fill_2
XFILLER_40_366 VPWR VGND sg13g2_fill_1
Xhold92 controller.const_data\[4\] VPWR VGND net419 sg13g2_dlygate4sd3_1
XFILLER_48_477 VPWR VGND sg13g2_decap_8
XFILLER_48_400 VPWR VGND sg13g2_decap_8
Xhold70 _0236_ VPWR VGND net397 sg13g2_dlygate4sd3_1
Xhold81 _0257_ VPWR VGND net408 sg13g2_dlygate4sd3_1
X_2830_ VGND VPWR _1054_ net569 _0215_ _0906_ sg13g2_a21oi_1
XANTENNA_1 VPWR VGND ui_in[0] sg13g2_antennanp
X_2761_ _0855_ net888 _1271_ VPWR VGND sg13g2_nand2_1
X_2692_ _0801_ _1063_ _0410_ VPWR VGND sg13g2_xnor2_1
X_1712_ _1063_ net879 VPWR VGND sg13g2_inv_2
X_1643_ VPWR _0994_ net847 VGND sg13g2_inv_1
X_3244_ net246 VGND VPWR net766 controller.inst_mem.mem_data\[59\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
Xfanout519 net522 net519 VPWR VGND sg13g2_buf_8
Xfanout508 net509 net508 VPWR VGND sg13g2_buf_2
X_3175_ net252 VGND VPWR net889 controller.counter2.counter_1\[6\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_1
XFILLER_39_466 VPWR VGND sg13g2_decap_8
X_2057_ net649 VPWR _0304_ VGND controller.inst_mem.mem_data\[126\] net596 sg13g2_o21ai_1
X_2126_ VGND VPWR _1137_ net546 _0079_ _0338_ sg13g2_a21oi_1
X_2959_ net662 VPWR _0971_ VGND controller.inst_mem.mem_data\[72\] net617 sg13g2_o21ai_1
XFILLER_45_414 VPWR VGND sg13g2_decap_8
XFILLER_13_377 VPWR VGND sg13g2_fill_1
XFILLER_36_447 VPWR VGND sg13g2_decap_8
XFILLER_0_281 VPWR VGND sg13g2_fill_1
X_2813_ net544 VPWR _0898_ VGND net909 net474 sg13g2_o21ai_1
X_2675_ net540 VPWR _0788_ VGND net928 net444 sg13g2_o21ai_1
X_2744_ net543 VPWR _0842_ VGND net911 net475 sg13g2_o21ai_1
X_3235__107 VPWR VGND net107 sg13g2_tiehi
X_3246__214 VPWR VGND net214 sg13g2_tiehi
X_3227_ net202 VGND VPWR _0250_ controller.inst_mem.mem_data\[42\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
X_3158_ net320 VGND VPWR net939 controller.counter2.counter_0\[5\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
XFILLER_42_428 VPWR VGND sg13g2_decap_8
X_3089_ net235 VGND VPWR _0112_ controller.inst_mem.mem_data\[193\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_2109_ net648 VPWR _0330_ VGND net771 net592 sg13g2_o21ai_1
X_3103__207 VPWR VGND net207 sg13g2_tiehi
Xhold392 _0181_ VPWR VGND net939 sg13g2_dlygate4sd3_1
Xhold381 controller.counter2.counter_0\[3\] VPWR VGND net928 sg13g2_dlygate4sd3_1
Xhold370 controller.output_controller.keep\[2\] VPWR VGND net917 sg13g2_dlygate4sd3_1
XFILLER_45_200 VPWR VGND sg13g2_fill_1
XFILLER_18_436 VPWR VGND sg13g2_fill_1
X_3160__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_26_93 VPWR VGND sg13g2_fill_1
X_3004__116 VPWR VGND net116 sg13g2_tiehi
X_2460_ VGND VPWR _0600_ _0601_ _0149_ _0602_ sg13g2_a21oi_1
XFILLER_9_189 VPWR VGND sg13g2_fill_2
X_2391_ _0533_ VPWR _0534_ VGND controller.inst_mem.mem_data\[54\] net491 sg13g2_o21ai_1
X_3012_ net100 VGND VPWR _0035_ controller.inst_mem.mem_data\[116\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_2658_ _0732_ _0768_ _0774_ VPWR VGND sg13g2_and2_1
X_2727_ VPWR VGND _0827_ net447 _0770_ net348 _0828_ net480 sg13g2_a221oi_1
X_2589_ _0709_ net7 _0581_ net483 VPWR VGND sg13g2_and3_1
XFILLER_2_365 VPWR VGND sg13g2_fill_2
XFILLER_33_203 VPWR VGND sg13g2_fill_1
X_1960_ _1305_ controller.alu_buffer.buffer\[22\] _1260_ VPWR VGND sg13g2_nand2_1
X_1891_ _1242_ _1238_ _1241_ net514 _1020_ VPWR VGND sg13g2_a22oi_1
X_2512_ net538 VPWR _0645_ VGND controller.alu_buffer.buffer\[10\] net460 sg13g2_o21ai_1
X_2443_ _0586_ net485 _0561_ _0581_ VPWR VGND sg13g2_and3_1
X_3056__301 VPWR VGND net301 sg13g2_tiehi
X_2374_ _0518_ net524 controller.extended_jump_target\[2\] net507 controller.inst_mem.mem_data\[58\]
+ VPWR VGND sg13g2_a22oi_1
X_2090_ VGND VPWR _1155_ net590 _0061_ _0320_ sg13g2_a21oi_1
X_2992_ net140 VGND VPWR _0015_ controller.inst_mem.mem_data\[96\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_1943_ _1284_ _1286_ _1283_ _1290_ VPWR VGND _1289_ sg13g2_nand4_1
X_1874_ _1225_ net534 net535 VPWR VGND sg13g2_nand2_1
X_2426_ _0566_ _0567_ _0565_ _0569_ VPWR VGND _0568_ sg13g2_nand4_1
XFILLER_37_394 VPWR VGND sg13g2_fill_1
X_2357_ _0503_ net637 VPWR VGND net6 sg13g2_nand2b_2
X_2288_ _0432_ _0433_ _0434_ VPWR VGND sg13g2_nor2_1
XFILLER_40_504 VPWR VGND sg13g2_decap_4
XFILLER_4_449 VPWR VGND sg13g2_fill_1
X_3260_ net302 VGND VPWR net367 controller.inst_mem.mem_data\[75\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
X_3191_ net188 VGND VPWR _0214_ controller.const_data\[6\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_38_147 VPWR VGND sg13g2_fill_2
X_2142_ VGND VPWR _1129_ net608 _0087_ _0346_ sg13g2_a21oi_1
X_2073_ net628 VPWR _0312_ VGND controller.inst_mem.mem_data\[134\] net557 sg13g2_o21ai_1
X_2211_ net645 VPWR _0381_ VGND net729 net582 sg13g2_o21ai_1
X_2975_ net648 VPWR _0979_ VGND net414 net594 sg13g2_o21ai_1
X_1926_ net901 controller.counter2.counter_1\[8\] controller.counter2.counter_1\[7\]
+ _1274_ VGND VPWR _1272_ sg13g2_nor4_2
X_1857_ VPWR _1208_ net370 VGND sg13g2_inv_1
X_3149__61 VPWR VGND net61 sg13g2_tiehi
X_1788_ VPWR _1139_ net867 VGND sg13g2_inv_1
X_2409_ VGND VPWR _0551_ _0552_ net517 _1005_ sg13g2_a21oi_2
Xhold93 _0213_ VPWR VGND net420 sg13g2_dlygate4sd3_1
XFILLER_48_456 VPWR VGND sg13g2_decap_8
Xhold82 controller.const_data\[18\] VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold71 controller.inst_mem.mem_data\[180\] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold60 _0033_ VPWR VGND net387 sg13g2_dlygate4sd3_1
XANTENNA_2 VPWR VGND ui_in[2] sg13g2_antennanp
X_2760_ VGND VPWR net476 _0853_ _0197_ _0854_ sg13g2_a21oi_1
X_2691_ VGND VPWR _0798_ _0799_ _0182_ _0800_ sg13g2_a21oi_1
X_1711_ VPWR _1062_ controller.counter2.counter_0\[10\] VGND sg13g2_inv_1
X_1642_ VPWR _0993_ net767 VGND sg13g2_inv_1
X_3243_ net262 VGND VPWR net427 controller.inst_mem.mem_data\[58\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
Xfanout509 _1220_ net509 VPWR VGND sg13g2_buf_8
X_3174_ net256 VGND VPWR _0197_ controller.counter2.counter_1\[5\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_1
XFILLER_39_445 VPWR VGND sg13g2_decap_8
X_2056_ VGND VPWR _1172_ net599 _0044_ _0303_ sg13g2_a21oi_1
X_2125_ net627 VPWR _0338_ VGND net402 net547 sg13g2_o21ai_1
X_2958_ VGND VPWR _0990_ net609 _0279_ _0970_ sg13g2_a21oi_1
X_3064__285 VPWR VGND net285 sg13g2_tiehi
X_1909_ _1235_ _1257_ _1260_ VPWR VGND sg13g2_nor2_2
X_2889_ net631 VPWR _0936_ VGND net869 net561 sg13g2_o21ai_1
X_3207__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_16_150 VPWR VGND sg13g2_fill_2
XFILLER_44_492 VPWR VGND sg13g2_decap_8
X_2743_ VGND VPWR net409 net451 _0841_ _0840_ sg13g2_a21oi_1
X_2812_ VGND VPWR net873 net450 _0897_ _0896_ sg13g2_a21oi_1
X_2674_ VPWR VGND net10 net446 _0774_ net838 _0787_ net479 sg13g2_a221oi_1
X_3157_ net324 VGND VPWR _0180_ controller.counter2.counter_0\[4\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_3226_ net210 VGND VPWR net723 controller.inst_mem.mem_data\[41\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_3088_ net237 VGND VPWR net395 controller.inst_mem.mem_data\[192\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_2108_ VGND VPWR _1146_ net594 _0070_ _0329_ sg13g2_a21oi_1
X_2039_ net655 VPWR _0295_ VGND controller.inst_mem.mem_data\[117\] net573 sg13g2_o21ai_1
XFILLER_22_164 VPWR VGND sg13g2_fill_2
Xhold382 _0179_ VPWR VGND net929 sg13g2_dlygate4sd3_1
Xhold360 controller.counter2.counter_1\[10\] VPWR VGND net907 sg13g2_dlygate4sd3_1
Xhold371 _0175_ VPWR VGND net918 sg13g2_dlygate4sd3_1
Xhold393 controller.output_controller.keep\[1\] VPWR VGND net940 sg13g2_dlygate4sd3_1
XFILLER_45_278 VPWR VGND sg13g2_fill_1
XFILLER_42_60 VPWR VGND sg13g2_fill_1
XFILLER_41_495 VPWR VGND sg13g2_decap_8
XFILLER_13_164 VPWR VGND sg13g2_fill_1
XFILLER_3_76 VPWR VGND sg13g2_fill_1
X_3011_ net102 VGND VPWR net764 controller.inst_mem.mem_data\[115\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_2390_ _0530_ _0531_ _0529_ _0533_ VPWR VGND _0532_ sg13g2_nand4_1
X_2726_ _0418_ net906 _0827_ VPWR VGND sg13g2_xor2_1
XFILLER_32_495 VPWR VGND sg13g2_decap_8
XFILLER_32_473 VPWR VGND sg13g2_decap_4
X_2657_ _0767_ VPWR _0773_ VGND _0732_ _0769_ sg13g2_o21ai_1
X_2588_ controller.alu_buffer.buffer\[22\] net485 _0561_ _0582_ _0708_ VPWR VGND sg13g2_and4_1
X_3209_ net63 VGND VPWR _0232_ controller.const_data\[24\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_42_226 VPWR VGND sg13g2_fill_2
XFILLER_10_156 VPWR VGND sg13g2_fill_2
Xhold190 controller.inst_mem.mem_data\[121\] VPWR VGND net737 sg13g2_dlygate4sd3_1
X_1890_ VPWR VGND controller.inst_mem.extended_word\[8\] _1240_ net523 controller.inst_mem.mem_data\[160\]
+ _1241_ net510 sg13g2_a221oi_1
X_2442_ _0585_ controller.alu_buffer.buffer\[7\] net472 VPWR VGND sg13g2_nand2_1
X_2511_ _0644_ net456 net933 net471 controller.alu_buffer.buffer\[9\] VPWR VGND sg13g2_a22oi_1
X_2373_ net488 VPWR _0517_ VGND net524 _0516_ sg13g2_o21ai_1
X_2709_ _0814_ net897 _0414_ VPWR VGND sg13g2_xnor2_1
X_1942_ controller.alu_buffer.buffer\[10\] controller.alu_buffer.buffer\[9\] controller.alu_buffer.buffer\[8\]
+ _1289_ VPWR VGND sg13g2_nor3_1
X_2991_ net142 VGND VPWR net802 controller.inst_mem.mem_data\[95\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_1873_ _1224_ net502 controller.inst_mem.mem_data\[183\] net506 controller.inst_mem.mem_data\[63\]
+ VPWR VGND sg13g2_a22oi_1
X_2356_ net6 net637 _0502_ VPWR VGND sg13g2_nor2b_2
X_2425_ _0568_ net495 controller.inst_mem.mem_data\[101\] net507 controller.inst_mem.mem_data\[77\]
+ VPWR VGND sg13g2_a22oi_1
X_2287_ controller.extended_cond.opcode\[1\] VPWR _0433_ VGND controller.extended_cond.opcode\[0\]
+ net3 sg13g2_o21ai_1
X_3074__265 VPWR VGND net265 sg13g2_tiehi
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
X_3190_ net192 VGND VPWR net420 controller.const_data\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2210_ VGND VPWR _1095_ net583 _0121_ _0380_ sg13g2_a21oi_1
X_2141_ net660 VPWR _0346_ VGND net336 net616 sg13g2_o21ai_1
X_2072_ VGND VPWR _1164_ net556 _0052_ _0311_ sg13g2_a21oi_1
X_1925_ VGND VPWR _1273_ _1272_ net932 sg13g2_or2_1
X_2974_ VGND VPWR _0982_ net595 _0287_ _0978_ sg13g2_a21oi_1
X_1787_ VPWR _1138_ net794 VGND sg13g2_inv_1
X_1856_ VPWR _1207_ net770 VGND sg13g2_inv_1
X_2408_ VGND VPWR controller.inst_mem.extended_word\[23\] net524 _0551_ _0550_ sg13g2_a21oi_1
X_2339_ VGND VPWR _0484_ _0485_ net515 _1024_ sg13g2_a21oi_2
X_3155__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_48_435 VPWR VGND sg13g2_decap_8
X_3163__300 VPWR VGND net300 sg13g2_tiehi
Xhold83 controller.const_data\[17\] VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold94 controller.inst_mem.mem_data\[97\] VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold72 _0100_ VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold61 controller.inst_mem.mem_data\[104\] VPWR VGND net388 sg13g2_dlygate4sd3_1
Xhold50 _0144_ VPWR VGND net377 sg13g2_dlygate4sd3_1
XFILLER_43_195 VPWR VGND sg13g2_fill_2
XANTENNA_3 VPWR VGND ui_in[3] sg13g2_antennanp
X_2690_ net539 VPWR _0800_ VGND net894 net444 sg13g2_o21ai_1
X_1710_ VPWR _1061_ net7 VGND sg13g2_inv_1
X_1641_ VPWR _0992_ net675 VGND sg13g2_inv_1
X_3173_ net260 VGND VPWR _0196_ controller.counter2.counter_1\[4\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_2
X_3242_ net278 VGND VPWR _0265_ controller.inst_mem.mem_data\[57\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_2124_ VGND VPWR _1138_ net546 _0078_ _0337_ sg13g2_a21oi_1
X_2055_ net652 VPWR _0303_ VGND net382 net599 sg13g2_o21ai_1
X_2957_ net656 VPWR _0970_ VGND net669 net609 sg13g2_o21ai_1
X_1839_ VPWR _1190_ net416 VGND sg13g2_inv_1
X_2888_ VGND VPWR _1025_ net582 _0244_ _0935_ sg13g2_a21oi_1
X_1908_ VGND VPWR _1248_ _1255_ _1259_ _1258_ sg13g2_a21oi_1
XFILLER_45_449 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_37_clk clknet_3_0__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_44_471 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_28_clk clknet_3_5__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
X_2742_ net454 _0839_ _0840_ VPWR VGND sg13g2_nor2_1
X_2811_ net450 _0895_ _0896_ VPWR VGND sg13g2_nor2_1
X_2673_ _0786_ net448 _0785_ VPWR VGND sg13g2_nand2b_1
X_3156_ net39 VGND VPWR net929 controller.counter2.counter_0\[3\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_3087_ net239 VGND VPWR net381 controller.inst_mem.mem_data\[191\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_19_clk clknet_3_7__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
X_2107_ net650 VPWR _0329_ VGND controller.inst_mem.mem_data\[151\] net593 sg13g2_o21ai_1
X_3225_ net218 VGND VPWR _0248_ controller.inst_mem.mem_data\[40\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
XFILLER_35_482 VPWR VGND sg13g2_decap_8
X_2038_ VGND VPWR _1181_ net565 _0035_ _0294_ sg13g2_a21oi_1
XFILLER_22_132 VPWR VGND sg13g2_fill_2
XFILLER_22_143 VPWR VGND sg13g2_fill_2
Xhold350 controller.counter2.counter_0\[11\] VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold372 controller.counter2.counter_0\[2\] VPWR VGND net919 sg13g2_dlygate4sd3_1
Xhold383 controller.counter2.counter_0\[1\] VPWR VGND net930 sg13g2_dlygate4sd3_1
Xhold361 _0202_ VPWR VGND net908 sg13g2_dlygate4sd3_1
Xhold394 _0174_ VPWR VGND net941 sg13g2_dlygate4sd3_1
XFILLER_41_474 VPWR VGND sg13g2_decap_8
X_3010_ net104 VGND VPWR net387 controller.inst_mem.mem_data\[114\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_3202__119 VPWR VGND net119 sg13g2_tiehi
X_2725_ _0825_ _0826_ _0190_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_2656_ _0766_ _0769_ net480 _0772_ VPWR VGND sg13g2_mux2_1
X_2587_ _0706_ net467 _0707_ VPWR VGND sg13g2_nor2b_1
X_3208_ net71 VGND VPWR _0231_ controller.const_data\[23\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3139_ net101 VGND VPWR net955 controller.alu_buffer.buffer\[13\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_27_279 VPWR VGND sg13g2_fill_1
Xhold180 _0263_ VPWR VGND net727 sg13g2_dlygate4sd3_1
Xfanout660 net662 net660 VPWR VGND sg13g2_buf_8
Xhold191 controller.inst_mem.mem_data\[174\] VPWR VGND net738 sg13g2_dlygate4sd3_1
XFILLER_26_290 VPWR VGND sg13g2_fill_1
X_3084__245 VPWR VGND net245 sg13g2_tiehi
X_2510_ VPWR VGND net467 net462 _0642_ controller.alu_buffer.buffer\[11\] _0643_ net482
+ sg13g2_a221oi_1
X_3019__86 VPWR VGND net86 sg13g2_tiehi
X_3034__56 VPWR VGND net56 sg13g2_tiehi
X_2441_ _0584_ net485 _0561_ _0582_ VPWR VGND sg13g2_and3_1
X_2372_ VGND VPWR net534 net535 _0516_ net531 sg13g2_a21oi_1
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_24_205 VPWR VGND sg13g2_fill_2
X_2708_ _0812_ _0813_ _0186_ VPWR VGND sg13g2_nor2_1
X_2639_ _0754_ VPWR _0755_ VGND net490 net489 sg13g2_o21ai_1
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_46_374 VPWR VGND sg13g2_decap_8
Xfanout490 _0422_ net490 VPWR VGND sg13g2_buf_2
X_1941_ VGND VPWR _1288_ _1287_ controller.alu_buffer.buffer\[8\] sg13g2_or2_1
X_2990_ net144 VGND VPWR net343 controller.inst_mem.mem_data\[94\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_1872_ net534 net531 _1223_ VPWR VGND net535 sg13g2_nand3b_1
XFILLER_36_0 VPWR VGND sg13g2_fill_1
X_2286_ net4 _0427_ _0432_ VPWR VGND sg13g2_nor2_1
X_2355_ _0477_ VPWR _0501_ VGND net486 _0500_ sg13g2_o21ai_1
X_2424_ VPWR VGND controller.inst_mem.mem_data\[149\] net517 net520 controller.inst_mem.mem_data\[125\]
+ _0567_ net499 sg13g2_a221oi_1
X_2140_ VGND VPWR _1130_ net608 _0086_ _0345_ sg13g2_a21oi_1
X_2071_ net628 VPWR _0311_ VGND net384 net556 sg13g2_o21ai_1
X_1924_ controller.counter2.counter_1\[6\] controller.counter2.counter_1\[5\] controller.counter2.counter_1\[4\]
+ _1270_ _1272_ VPWR VGND sg13g2_or4_1
X_2973_ net650 VPWR _0978_ VGND net691 net595 sg13g2_o21ai_1
X_1855_ VPWR _1206_ net423 VGND sg13g2_inv_1
X_1786_ VPWR _1137_ net871 VGND sg13g2_inv_1
X_2269_ VGND VPWR _0415_ _0414_ net897 sg13g2_or2_1
X_3110__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_25_300 VPWR VGND sg13g2_fill_2
X_2407_ _0548_ _0549_ _0547_ _0550_ VPWR VGND sg13g2_nand3_1
X_2338_ _0484_ _1280_ _0483_ VPWR VGND sg13g2_nand2_1
XFILLER_40_347 VPWR VGND sg13g2_fill_1
XFILLER_48_414 VPWR VGND sg13g2_decap_8
Xhold40 _0283_ VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold73 controller.inst_mem.mem_data\[194\] VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold95 _0017_ VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold62 _0024_ VPWR VGND net389 sg13g2_dlygate4sd3_1
Xhold51 controller.inst_mem.mem_data\[183\] VPWR VGND net378 sg13g2_dlygate4sd3_1
Xhold84 controller.inst_mem.mem_data\[139\] VPWR VGND net411 sg13g2_dlygate4sd3_1
XFILLER_16_366 VPWR VGND sg13g2_fill_1
XFILLER_31_358 VPWR VGND sg13g2_fill_1
XANTENNA_4 VPWR VGND ui_in[5] sg13g2_antennanp
X_1640_ VPWR _0991_ net857 VGND sg13g2_inv_1
XFILLER_6_33 VPWR VGND sg13g2_fill_2
X_3172_ net264 VGND VPWR net891 controller.counter2.counter_1\[3\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_1
X_2123_ net627 VPWR _0337_ VGND controller.inst_mem.mem_data\[159\] net546 sg13g2_o21ai_1
X_3241_ net294 VGND VPWR _0264_ controller.inst_mem.mem_data\[56\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_2054_ VGND VPWR _1173_ net602 _0043_ _0302_ sg13g2_a21oi_1
X_2956_ VGND VPWR _0991_ net606 _0278_ _0969_ sg13g2_a21oi_1
X_1838_ VPWR _1189_ net775 VGND sg13g2_inv_1
X_2887_ net645 VPWR _0935_ VGND controller.inst_mem.mem_data\[36\] net561 sg13g2_o21ai_1
X_1907_ _1236_ _1257_ _1258_ VPWR VGND sg13g2_nor2_2
X_1769_ VPWR _1120_ net850 VGND sg13g2_inv_1
XFILLER_45_428 VPWR VGND sg13g2_decap_8
XFILLER_40_122 VPWR VGND sg13g2_fill_1
X_3043__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_13_314 VPWR VGND sg13g2_fill_2
XFILLER_44_450 VPWR VGND sg13g2_decap_8
X_2672_ _0785_ net928 _0406_ VPWR VGND sg13g2_xnor2_1
X_2741_ _1269_ _0838_ _0839_ VPWR VGND sg13g2_nor2b_1
X_2810_ VGND VPWR net909 _0890_ _0895_ _1279_ sg13g2_a21oi_1
X_3094__225 VPWR VGND net225 sg13g2_tiehi
X_3224_ net226 VGND VPWR _0247_ controller.inst_mem.mem_data\[39\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
.ends

