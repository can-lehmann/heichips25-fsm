module heichips25_can_lehmann_fsm (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire clknet_leaf_0_clk;
 wire \controller.alu_buffer.buffer[0] ;
 wire \controller.alu_buffer.buffer[10] ;
 wire \controller.alu_buffer.buffer[11] ;
 wire \controller.alu_buffer.buffer[12] ;
 wire \controller.alu_buffer.buffer[13] ;
 wire \controller.alu_buffer.buffer[14] ;
 wire \controller.alu_buffer.buffer[15] ;
 wire \controller.alu_buffer.buffer[16] ;
 wire \controller.alu_buffer.buffer[17] ;
 wire \controller.alu_buffer.buffer[18] ;
 wire \controller.alu_buffer.buffer[19] ;
 wire \controller.alu_buffer.buffer[1] ;
 wire \controller.alu_buffer.buffer[20] ;
 wire \controller.alu_buffer.buffer[21] ;
 wire \controller.alu_buffer.buffer[22] ;
 wire \controller.alu_buffer.buffer[23] ;
 wire \controller.alu_buffer.buffer[2] ;
 wire \controller.alu_buffer.buffer[3] ;
 wire \controller.alu_buffer.buffer[4] ;
 wire \controller.alu_buffer.buffer[5] ;
 wire \controller.alu_buffer.buffer[6] ;
 wire \controller.alu_buffer.buffer[7] ;
 wire \controller.alu_buffer.buffer[8] ;
 wire \controller.alu_buffer.buffer[9] ;
 wire \controller.const_data[0] ;
 wire \controller.const_data[10] ;
 wire \controller.const_data[11] ;
 wire \controller.const_data[12] ;
 wire \controller.const_data[13] ;
 wire \controller.const_data[14] ;
 wire \controller.const_data[15] ;
 wire \controller.const_data[16] ;
 wire \controller.const_data[17] ;
 wire \controller.const_data[18] ;
 wire \controller.const_data[19] ;
 wire \controller.const_data[1] ;
 wire \controller.const_data[20] ;
 wire \controller.const_data[21] ;
 wire \controller.const_data[22] ;
 wire \controller.const_data[23] ;
 wire \controller.const_data[24] ;
 wire \controller.const_data[25] ;
 wire \controller.const_data[26] ;
 wire \controller.const_data[27] ;
 wire \controller.const_data[28] ;
 wire \controller.const_data[29] ;
 wire \controller.const_data[2] ;
 wire \controller.const_data[30] ;
 wire \controller.const_data[31] ;
 wire \controller.const_data[3] ;
 wire \controller.const_data[4] ;
 wire \controller.const_data[5] ;
 wire \controller.const_data[6] ;
 wire \controller.const_data[7] ;
 wire \controller.const_data[8] ;
 wire \controller.const_data[9] ;
 wire \controller.counter2.counter_0[0] ;
 wire \controller.counter2.counter_0[10] ;
 wire \controller.counter2.counter_0[11] ;
 wire \controller.counter2.counter_0[12] ;
 wire \controller.counter2.counter_0[13] ;
 wire \controller.counter2.counter_0[14] ;
 wire \controller.counter2.counter_0[15] ;
 wire \controller.counter2.counter_0[1] ;
 wire \controller.counter2.counter_0[2] ;
 wire \controller.counter2.counter_0[3] ;
 wire \controller.counter2.counter_0[4] ;
 wire \controller.counter2.counter_0[5] ;
 wire \controller.counter2.counter_0[6] ;
 wire \controller.counter2.counter_0[7] ;
 wire \controller.counter2.counter_0[8] ;
 wire \controller.counter2.counter_0[9] ;
 wire \controller.counter2.counter_1[0] ;
 wire \controller.counter2.counter_1[10] ;
 wire \controller.counter2.counter_1[11] ;
 wire \controller.counter2.counter_1[12] ;
 wire \controller.counter2.counter_1[13] ;
 wire \controller.counter2.counter_1[14] ;
 wire \controller.counter2.counter_1[15] ;
 wire \controller.counter2.counter_1[1] ;
 wire \controller.counter2.counter_1[2] ;
 wire \controller.counter2.counter_1[3] ;
 wire \controller.counter2.counter_1[4] ;
 wire \controller.counter2.counter_1[5] ;
 wire \controller.counter2.counter_1[6] ;
 wire \controller.counter2.counter_1[7] ;
 wire \controller.counter2.counter_1[8] ;
 wire \controller.counter2.counter_1[9] ;
 wire \controller.extended_cond.opcode[0] ;
 wire \controller.extended_cond.opcode[1] ;
 wire \controller.extended_cond.opcode[2] ;
 wire \controller.extended_jump_target[0] ;
 wire \controller.extended_jump_target[1] ;
 wire \controller.extended_jump_target[2] ;
 wire \controller.extended_state[0] ;
 wire \controller.extended_state[1] ;
 wire \controller.extended_state[2] ;
 wire \controller.extended_then_action[0] ;
 wire \controller.extended_then_action[1] ;
 wire \controller.extended_then_action[2] ;
 wire \controller.extended_then_action[3] ;
 wire \controller.extended_then_action[4] ;
 wire \controller.extended_then_action[5] ;
 wire \controller.inst_mem.addr[0] ;
 wire \controller.inst_mem.addr[1] ;
 wire \controller.inst_mem.addr[2] ;
 wire \controller.inst_mem.extended_word[18] ;
 wire \controller.inst_mem.extended_word[19] ;
 wire \controller.inst_mem.extended_word[20] ;
 wire \controller.inst_mem.extended_word[21] ;
 wire \controller.inst_mem.extended_word[22] ;
 wire \controller.inst_mem.extended_word[23] ;
 wire \controller.inst_mem.extended_word[3] ;
 wire \controller.inst_mem.extended_word[4] ;
 wire \controller.inst_mem.extended_word[5] ;
 wire \controller.inst_mem.extended_word[6] ;
 wire \controller.inst_mem.extended_word[7] ;
 wire \controller.inst_mem.extended_word[8] ;
 wire \controller.inst_mem.mem_data[100] ;
 wire \controller.inst_mem.mem_data[101] ;
 wire \controller.inst_mem.mem_data[102] ;
 wire \controller.inst_mem.mem_data[103] ;
 wire \controller.inst_mem.mem_data[104] ;
 wire \controller.inst_mem.mem_data[105] ;
 wire \controller.inst_mem.mem_data[106] ;
 wire \controller.inst_mem.mem_data[107] ;
 wire \controller.inst_mem.mem_data[108] ;
 wire \controller.inst_mem.mem_data[109] ;
 wire \controller.inst_mem.mem_data[110] ;
 wire \controller.inst_mem.mem_data[111] ;
 wire \controller.inst_mem.mem_data[112] ;
 wire \controller.inst_mem.mem_data[113] ;
 wire \controller.inst_mem.mem_data[114] ;
 wire \controller.inst_mem.mem_data[115] ;
 wire \controller.inst_mem.mem_data[116] ;
 wire \controller.inst_mem.mem_data[117] ;
 wire \controller.inst_mem.mem_data[118] ;
 wire \controller.inst_mem.mem_data[119] ;
 wire \controller.inst_mem.mem_data[120] ;
 wire \controller.inst_mem.mem_data[121] ;
 wire \controller.inst_mem.mem_data[122] ;
 wire \controller.inst_mem.mem_data[123] ;
 wire \controller.inst_mem.mem_data[124] ;
 wire \controller.inst_mem.mem_data[125] ;
 wire \controller.inst_mem.mem_data[126] ;
 wire \controller.inst_mem.mem_data[127] ;
 wire \controller.inst_mem.mem_data[128] ;
 wire \controller.inst_mem.mem_data[129] ;
 wire \controller.inst_mem.mem_data[130] ;
 wire \controller.inst_mem.mem_data[131] ;
 wire \controller.inst_mem.mem_data[132] ;
 wire \controller.inst_mem.mem_data[133] ;
 wire \controller.inst_mem.mem_data[134] ;
 wire \controller.inst_mem.mem_data[135] ;
 wire \controller.inst_mem.mem_data[136] ;
 wire \controller.inst_mem.mem_data[137] ;
 wire \controller.inst_mem.mem_data[138] ;
 wire \controller.inst_mem.mem_data[139] ;
 wire \controller.inst_mem.mem_data[140] ;
 wire \controller.inst_mem.mem_data[141] ;
 wire \controller.inst_mem.mem_data[142] ;
 wire \controller.inst_mem.mem_data[143] ;
 wire \controller.inst_mem.mem_data[144] ;
 wire \controller.inst_mem.mem_data[145] ;
 wire \controller.inst_mem.mem_data[146] ;
 wire \controller.inst_mem.mem_data[147] ;
 wire \controller.inst_mem.mem_data[148] ;
 wire \controller.inst_mem.mem_data[149] ;
 wire \controller.inst_mem.mem_data[150] ;
 wire \controller.inst_mem.mem_data[151] ;
 wire \controller.inst_mem.mem_data[152] ;
 wire \controller.inst_mem.mem_data[153] ;
 wire \controller.inst_mem.mem_data[154] ;
 wire \controller.inst_mem.mem_data[155] ;
 wire \controller.inst_mem.mem_data[156] ;
 wire \controller.inst_mem.mem_data[157] ;
 wire \controller.inst_mem.mem_data[158] ;
 wire \controller.inst_mem.mem_data[159] ;
 wire \controller.inst_mem.mem_data[160] ;
 wire \controller.inst_mem.mem_data[161] ;
 wire \controller.inst_mem.mem_data[162] ;
 wire \controller.inst_mem.mem_data[163] ;
 wire \controller.inst_mem.mem_data[164] ;
 wire \controller.inst_mem.mem_data[165] ;
 wire \controller.inst_mem.mem_data[166] ;
 wire \controller.inst_mem.mem_data[167] ;
 wire \controller.inst_mem.mem_data[168] ;
 wire \controller.inst_mem.mem_data[169] ;
 wire \controller.inst_mem.mem_data[170] ;
 wire \controller.inst_mem.mem_data[171] ;
 wire \controller.inst_mem.mem_data[172] ;
 wire \controller.inst_mem.mem_data[173] ;
 wire \controller.inst_mem.mem_data[174] ;
 wire \controller.inst_mem.mem_data[175] ;
 wire \controller.inst_mem.mem_data[176] ;
 wire \controller.inst_mem.mem_data[177] ;
 wire \controller.inst_mem.mem_data[178] ;
 wire \controller.inst_mem.mem_data[179] ;
 wire \controller.inst_mem.mem_data[180] ;
 wire \controller.inst_mem.mem_data[181] ;
 wire \controller.inst_mem.mem_data[182] ;
 wire \controller.inst_mem.mem_data[183] ;
 wire \controller.inst_mem.mem_data[184] ;
 wire \controller.inst_mem.mem_data[185] ;
 wire \controller.inst_mem.mem_data[186] ;
 wire \controller.inst_mem.mem_data[187] ;
 wire \controller.inst_mem.mem_data[188] ;
 wire \controller.inst_mem.mem_data[189] ;
 wire \controller.inst_mem.mem_data[190] ;
 wire \controller.inst_mem.mem_data[191] ;
 wire \controller.inst_mem.mem_data[192] ;
 wire \controller.inst_mem.mem_data[193] ;
 wire \controller.inst_mem.mem_data[194] ;
 wire \controller.inst_mem.mem_data[195] ;
 wire \controller.inst_mem.mem_data[196] ;
 wire \controller.inst_mem.mem_data[197] ;
 wire \controller.inst_mem.mem_data[198] ;
 wire \controller.inst_mem.mem_data[199] ;
 wire \controller.inst_mem.mem_data[32] ;
 wire \controller.inst_mem.mem_data[33] ;
 wire \controller.inst_mem.mem_data[34] ;
 wire \controller.inst_mem.mem_data[35] ;
 wire \controller.inst_mem.mem_data[36] ;
 wire \controller.inst_mem.mem_data[37] ;
 wire \controller.inst_mem.mem_data[38] ;
 wire \controller.inst_mem.mem_data[39] ;
 wire \controller.inst_mem.mem_data[40] ;
 wire \controller.inst_mem.mem_data[41] ;
 wire \controller.inst_mem.mem_data[42] ;
 wire \controller.inst_mem.mem_data[43] ;
 wire \controller.inst_mem.mem_data[44] ;
 wire \controller.inst_mem.mem_data[45] ;
 wire \controller.inst_mem.mem_data[46] ;
 wire \controller.inst_mem.mem_data[47] ;
 wire \controller.inst_mem.mem_data[48] ;
 wire \controller.inst_mem.mem_data[49] ;
 wire \controller.inst_mem.mem_data[50] ;
 wire \controller.inst_mem.mem_data[51] ;
 wire \controller.inst_mem.mem_data[52] ;
 wire \controller.inst_mem.mem_data[53] ;
 wire \controller.inst_mem.mem_data[54] ;
 wire \controller.inst_mem.mem_data[55] ;
 wire \controller.inst_mem.mem_data[56] ;
 wire \controller.inst_mem.mem_data[57] ;
 wire \controller.inst_mem.mem_data[58] ;
 wire \controller.inst_mem.mem_data[59] ;
 wire \controller.inst_mem.mem_data[60] ;
 wire \controller.inst_mem.mem_data[61] ;
 wire \controller.inst_mem.mem_data[62] ;
 wire \controller.inst_mem.mem_data[63] ;
 wire \controller.inst_mem.mem_data[64] ;
 wire \controller.inst_mem.mem_data[65] ;
 wire \controller.inst_mem.mem_data[66] ;
 wire \controller.inst_mem.mem_data[67] ;
 wire \controller.inst_mem.mem_data[68] ;
 wire \controller.inst_mem.mem_data[69] ;
 wire \controller.inst_mem.mem_data[70] ;
 wire \controller.inst_mem.mem_data[71] ;
 wire \controller.inst_mem.mem_data[72] ;
 wire \controller.inst_mem.mem_data[73] ;
 wire \controller.inst_mem.mem_data[74] ;
 wire \controller.inst_mem.mem_data[75] ;
 wire \controller.inst_mem.mem_data[76] ;
 wire \controller.inst_mem.mem_data[77] ;
 wire \controller.inst_mem.mem_data[78] ;
 wire \controller.inst_mem.mem_data[79] ;
 wire \controller.inst_mem.mem_data[80] ;
 wire \controller.inst_mem.mem_data[81] ;
 wire \controller.inst_mem.mem_data[82] ;
 wire \controller.inst_mem.mem_data[83] ;
 wire \controller.inst_mem.mem_data[84] ;
 wire \controller.inst_mem.mem_data[85] ;
 wire \controller.inst_mem.mem_data[86] ;
 wire \controller.inst_mem.mem_data[87] ;
 wire \controller.inst_mem.mem_data[88] ;
 wire \controller.inst_mem.mem_data[89] ;
 wire \controller.inst_mem.mem_data[90] ;
 wire \controller.inst_mem.mem_data[91] ;
 wire \controller.inst_mem.mem_data[92] ;
 wire \controller.inst_mem.mem_data[93] ;
 wire \controller.inst_mem.mem_data[94] ;
 wire \controller.inst_mem.mem_data[95] ;
 wire \controller.inst_mem.mem_data[96] ;
 wire \controller.inst_mem.mem_data[97] ;
 wire \controller.inst_mem.mem_data[98] ;
 wire \controller.inst_mem.mem_data[99] ;
 wire \controller.output_controller.keep[0] ;
 wire \controller.output_controller.keep[1] ;
 wire \controller.output_controller.keep[2] ;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net23;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;

 sg13g2_inv_1 _1629_ (.VDD(VPWR),
    .Y(_0980_),
    .A(net414),
    .VSS(VGND));
 sg13g2_inv_1 _1630_ (.VDD(VPWR),
    .Y(_0981_),
    .A(net691),
    .VSS(VGND));
 sg13g2_inv_1 _1631_ (.VDD(VPWR),
    .Y(_0982_),
    .A(net874),
    .VSS(VGND));
 sg13g2_inv_1 _1632_ (.VDD(VPWR),
    .Y(_0983_),
    .A(net826),
    .VSS(VGND));
 sg13g2_inv_1 _1633_ (.VDD(VPWR),
    .Y(_0984_),
    .A(net835),
    .VSS(VGND));
 sg13g2_inv_1 _1634_ (.VDD(VPWR),
    .Y(_0985_),
    .A(net792),
    .VSS(VGND));
 sg13g2_inv_1 _1635_ (.VDD(VPWR),
    .Y(_0986_),
    .A(net366),
    .VSS(VGND));
 sg13g2_inv_1 _1636_ (.VDD(VPWR),
    .Y(_0987_),
    .A(net346),
    .VSS(VGND));
 sg13g2_inv_1 _1637_ (.VDD(VPWR),
    .Y(_0988_),
    .A(net734),
    .VSS(VGND));
 sg13g2_inv_1 _1638_ (.VDD(VPWR),
    .Y(_0989_),
    .A(net669),
    .VSS(VGND));
 sg13g2_inv_1 _1639_ (.VDD(VPWR),
    .Y(_0990_),
    .A(net803),
    .VSS(VGND));
 sg13g2_inv_1 _1640_ (.VDD(VPWR),
    .Y(_0991_),
    .A(net857),
    .VSS(VGND));
 sg13g2_inv_1 _1641_ (.VDD(VPWR),
    .Y(_0992_),
    .A(net675),
    .VSS(VGND));
 sg13g2_inv_1 _1642_ (.VDD(VPWR),
    .Y(_0993_),
    .A(net767),
    .VSS(VGND));
 sg13g2_inv_1 _1643_ (.VDD(VPWR),
    .Y(_0994_),
    .A(net847),
    .VSS(VGND));
 sg13g2_inv_1 _1644_ (.VDD(VPWR),
    .Y(_0995_),
    .A(net374),
    .VSS(VGND));
 sg13g2_inv_1 _1645_ (.VDD(VPWR),
    .Y(_0996_),
    .A(net328),
    .VSS(VGND));
 sg13g2_inv_1 _1646_ (.VDD(VPWR),
    .Y(_0997_),
    .A(net862),
    .VSS(VGND));
 sg13g2_inv_1 _1647_ (.VDD(VPWR),
    .Y(_0998_),
    .A(net758),
    .VSS(VGND));
 sg13g2_inv_1 _1648_ (.VDD(VPWR),
    .Y(_0999_),
    .A(net864),
    .VSS(VGND));
 sg13g2_inv_1 _1649_ (.VDD(VPWR),
    .Y(_1000_),
    .A(net807),
    .VSS(VGND));
 sg13g2_inv_1 _1650_ (.VDD(VPWR),
    .Y(_1001_),
    .A(net809),
    .VSS(VGND));
 sg13g2_inv_1 _1651_ (.VDD(VPWR),
    .Y(_1002_),
    .A(net765),
    .VSS(VGND));
 sg13g2_inv_1 _1652_ (.VDD(VPWR),
    .Y(_1003_),
    .A(net426),
    .VSS(VGND));
 sg13g2_inv_1 _1653_ (.VDD(VPWR),
    .Y(_1004_),
    .A(net804),
    .VSS(VGND));
 sg13g2_inv_1 _1654_ (.VDD(VPWR),
    .Y(_1005_),
    .A(net872),
    .VSS(VGND));
 sg13g2_inv_1 _1655_ (.VDD(VPWR),
    .Y(_1006_),
    .A(net726),
    .VSS(VGND));
 sg13g2_inv_1 _1656_ (.VDD(VPWR),
    .Y(_1007_),
    .A(net812),
    .VSS(VGND));
 sg13g2_inv_1 _1657_ (.VDD(VPWR),
    .Y(_1008_),
    .A(net786),
    .VSS(VGND));
 sg13g2_inv_1 _1658_ (.VDD(VPWR),
    .Y(_1009_),
    .A(net432),
    .VSS(VGND));
 sg13g2_inv_1 _1659_ (.VDD(VPWR),
    .Y(_1010_),
    .A(net434),
    .VSS(VGND));
 sg13g2_inv_1 _1660_ (.VDD(VPWR),
    .Y(_1011_),
    .A(net852),
    .VSS(VGND));
 sg13g2_inv_1 _1661_ (.VDD(VPWR),
    .Y(_1012_),
    .A(net407),
    .VSS(VGND));
 sg13g2_inv_1 _1662_ (.VDD(VPWR),
    .Y(_1013_),
    .A(net413),
    .VSS(VGND));
 sg13g2_inv_1 _1663_ (.VDD(VPWR),
    .Y(_1014_),
    .A(net750),
    .VSS(VGND));
 sg13g2_inv_1 _1664_ (.VDD(VPWR),
    .Y(_1015_),
    .A(net664),
    .VSS(VGND));
 sg13g2_inv_1 _1665_ (.VDD(VPWR),
    .Y(_1016_),
    .A(net693),
    .VSS(VGND));
 sg13g2_inv_1 _1666_ (.VDD(VPWR),
    .Y(_1017_),
    .A(net853),
    .VSS(VGND));
 sg13g2_inv_1 _1667_ (.VDD(VPWR),
    .Y(_1018_),
    .A(net740),
    .VSS(VGND));
 sg13g2_inv_1 _1668_ (.VDD(VPWR),
    .Y(_1019_),
    .A(net856),
    .VSS(VGND));
 sg13g2_inv_1 _1669_ (.VDD(VPWR),
    .Y(_1020_),
    .A(net722),
    .VSS(VGND));
 sg13g2_inv_1 _1670_ (.VDD(VPWR),
    .Y(_1021_),
    .A(net799),
    .VSS(VGND));
 sg13g2_inv_1 _1671_ (.VDD(VPWR),
    .Y(_1022_),
    .A(net877),
    .VSS(VGND));
 sg13g2_inv_1 _1672_ (.VDD(VPWR),
    .Y(_1023_),
    .A(net869),
    .VSS(VGND));
 sg13g2_inv_2 _1673_ (.Y(_1024_),
    .A(net876),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1674_ (.VDD(VPWR),
    .Y(_1025_),
    .A(net748),
    .VSS(VGND));
 sg13g2_inv_1 _1675_ (.VDD(VPWR),
    .Y(_1026_),
    .A(net800),
    .VSS(VGND));
 sg13g2_inv_1 _1676_ (.VDD(VPWR),
    .Y(_1027_),
    .A(net720),
    .VSS(VGND));
 sg13g2_inv_1 _1677_ (.VDD(VPWR),
    .Y(_1028_),
    .A(net777),
    .VSS(VGND));
 sg13g2_inv_1 _1678_ (.VDD(VPWR),
    .Y(_1029_),
    .A(net873),
    .VSS(VGND));
 sg13g2_inv_1 _1679_ (.VDD(VPWR),
    .Y(_1030_),
    .A(net689),
    .VSS(VGND));
 sg13g2_inv_1 _1680_ (.VDD(VPWR),
    .Y(_1031_),
    .A(net440),
    .VSS(VGND));
 sg13g2_inv_1 _1681_ (.VDD(VPWR),
    .Y(_1032_),
    .A(net822),
    .VSS(VGND));
 sg13g2_inv_1 _1682_ (.VDD(VPWR),
    .Y(_1033_),
    .A(net396),
    .VSS(VGND));
 sg13g2_inv_1 _1683_ (.VDD(VPWR),
    .Y(_1034_),
    .A(net818),
    .VSS(VGND));
 sg13g2_inv_1 _1684_ (.VDD(VPWR),
    .Y(_1035_),
    .A(net687),
    .VSS(VGND));
 sg13g2_inv_1 _1685_ (.VDD(VPWR),
    .Y(_1036_),
    .A(net811),
    .VSS(VGND));
 sg13g2_inv_1 _1686_ (.VDD(VPWR),
    .Y(_1037_),
    .A(net820),
    .VSS(VGND));
 sg13g2_inv_1 _1687_ (.VDD(VPWR),
    .Y(_1038_),
    .A(net840),
    .VSS(VGND));
 sg13g2_inv_1 _1688_ (.VDD(VPWR),
    .Y(_1039_),
    .A(net718),
    .VSS(VGND));
 sg13g2_inv_1 _1689_ (.VDD(VPWR),
    .Y(_1040_),
    .A(net736),
    .VSS(VGND));
 sg13g2_inv_1 _1690_ (.VDD(VPWR),
    .Y(_1041_),
    .A(net344),
    .VSS(VGND));
 sg13g2_inv_1 _1691_ (.VDD(VPWR),
    .Y(_1042_),
    .A(net409),
    .VSS(VGND));
 sg13g2_inv_1 _1692_ (.VDD(VPWR),
    .Y(_1043_),
    .A(net410),
    .VSS(VGND));
 sg13g2_inv_1 _1693_ (.VDD(VPWR),
    .Y(_1044_),
    .A(net418),
    .VSS(VGND));
 sg13g2_inv_1 _1694_ (.VDD(VPWR),
    .Y(_1045_),
    .A(net348),
    .VSS(VGND));
 sg13g2_inv_1 _1695_ (.VDD(VPWR),
    .Y(_1046_),
    .A(net694),
    .VSS(VGND));
 sg13g2_inv_1 _1696_ (.VDD(VPWR),
    .Y(_1047_),
    .A(net707),
    .VSS(VGND));
 sg13g2_inv_1 _1697_ (.VDD(VPWR),
    .Y(_1048_),
    .A(net372),
    .VSS(VGND));
 sg13g2_inv_1 _1698_ (.VDD(VPWR),
    .Y(_1049_),
    .A(net681),
    .VSS(VGND));
 sg13g2_inv_1 _1699_ (.VDD(VPWR),
    .Y(_1050_),
    .A(net713),
    .VSS(VGND));
 sg13g2_inv_1 _1700_ (.VDD(VPWR),
    .Y(_1051_),
    .A(net390),
    .VSS(VGND));
 sg13g2_inv_1 _1701_ (.VDD(VPWR),
    .Y(_1052_),
    .A(net788),
    .VSS(VGND));
 sg13g2_inv_1 _1702_ (.VDD(VPWR),
    .Y(_1053_),
    .A(net824),
    .VSS(VGND));
 sg13g2_inv_1 _1703_ (.VDD(VPWR),
    .Y(_1054_),
    .A(net715),
    .VSS(VGND));
 sg13g2_inv_1 _1704_ (.VDD(VPWR),
    .Y(_1055_),
    .A(net774),
    .VSS(VGND));
 sg13g2_inv_1 _1705_ (.VDD(VPWR),
    .Y(_1056_),
    .A(net419),
    .VSS(VGND));
 sg13g2_inv_1 _1706_ (.VDD(VPWR),
    .Y(_1057_),
    .A(net838),
    .VSS(VGND));
 sg13g2_inv_1 _1707_ (.VDD(VPWR),
    .Y(_1058_),
    .A(net832),
    .VSS(VGND));
 sg13g2_inv_1 _1708_ (.VDD(VPWR),
    .Y(_1059_),
    .A(net695),
    .VSS(VGND));
 sg13g2_inv_1 _1709_ (.VDD(VPWR),
    .Y(_1060_),
    .A(net671),
    .VSS(VGND));
 sg13g2_inv_1 _1710_ (.VDD(VPWR),
    .Y(_1061_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _1711_ (.VDD(VPWR),
    .Y(_1062_),
    .A(\controller.counter2.counter_0[10] ),
    .VSS(VGND));
 sg13g2_inv_2 _1712_ (.Y(_1063_),
    .A(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _1713_ (.Y(_1064_),
    .A(net922),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1714_ (.VDD(VPWR),
    .Y(_1065_),
    .A(net963),
    .VSS(VGND));
 sg13g2_inv_1 _1715_ (.VDD(VPWR),
    .Y(_1066_),
    .A(\controller.alu_buffer.buffer[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _1716_ (.VDD(VPWR),
    .Y(_1067_),
    .A(net971),
    .VSS(VGND));
 sg13g2_inv_2 _1717_ (.Y(_1068_),
    .A(net531),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1718_ (.VDD(VPWR),
    .Y(_1069_),
    .A(net533),
    .VSS(VGND));
 sg13g2_inv_1 _1719_ (.VDD(VPWR),
    .Y(_1070_),
    .A(net535),
    .VSS(VGND));
 sg13g2_inv_1 _1720_ (.VDD(VPWR),
    .Y(_1071_),
    .A(net751),
    .VSS(VGND));
 sg13g2_inv_1 _1721_ (.VDD(VPWR),
    .Y(_1072_),
    .A(net376),
    .VSS(VGND));
 sg13g2_inv_1 _1722_ (.VDD(VPWR),
    .Y(_1073_),
    .A(net783),
    .VSS(VGND));
 sg13g2_inv_1 _1723_ (.VDD(VPWR),
    .Y(_1074_),
    .A(net353),
    .VSS(VGND));
 sg13g2_inv_1 _1724_ (.VDD(VPWR),
    .Y(_1075_),
    .A(net683),
    .VSS(VGND));
 sg13g2_inv_1 _1725_ (.VDD(VPWR),
    .Y(_1076_),
    .A(net403),
    .VSS(VGND));
 sg13g2_inv_1 _1726_ (.VDD(VPWR),
    .Y(_1077_),
    .A(net392),
    .VSS(VGND));
 sg13g2_inv_1 _1727_ (.VDD(VPWR),
    .Y(_1078_),
    .A(net364),
    .VSS(VGND));
 sg13g2_inv_2 _1728_ (.Y(_1079_),
    .A(net878),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1729_ (.VDD(VPWR),
    .Y(_1080_),
    .A(net881),
    .VSS(VGND));
 sg13g2_inv_1 _1730_ (.VDD(VPWR),
    .Y(_1081_),
    .A(net882),
    .VSS(VGND));
 sg13g2_inv_1 _1731_ (.VDD(VPWR),
    .Y(_1082_),
    .A(net685),
    .VSS(VGND));
 sg13g2_inv_1 _1732_ (.VDD(VPWR),
    .Y(_1083_),
    .A(net728),
    .VSS(VGND));
 sg13g2_inv_1 _1733_ (.VDD(VPWR),
    .Y(_1084_),
    .A(net858),
    .VSS(VGND));
 sg13g2_inv_1 _1734_ (.VDD(VPWR),
    .Y(_1085_),
    .A(net885),
    .VSS(VGND));
 sg13g2_inv_1 _1735_ (.VDD(VPWR),
    .Y(_1086_),
    .A(net943),
    .VSS(VGND));
 sg13g2_inv_1 _1736_ (.VDD(VPWR),
    .Y(_1087_),
    .A(net936),
    .VSS(VGND));
 sg13g2_inv_1 _1737_ (.VDD(VPWR),
    .Y(_1088_),
    .A(net761),
    .VSS(VGND));
 sg13g2_inv_1 _1738_ (.VDD(VPWR),
    .Y(_1089_),
    .A(net782),
    .VSS(VGND));
 sg13g2_inv_1 _1739_ (.VDD(VPWR),
    .Y(_1090_),
    .A(net701),
    .VSS(VGND));
 sg13g2_inv_1 _1740_ (.VDD(VPWR),
    .Y(_1091_),
    .A(net710),
    .VSS(VGND));
 sg13g2_inv_1 _1741_ (.VDD(VPWR),
    .Y(_1092_),
    .A(net334),
    .VSS(VGND));
 sg13g2_inv_1 _1742_ (.VDD(VPWR),
    .Y(_1093_),
    .A(net729),
    .VSS(VGND));
 sg13g2_inv_1 _1743_ (.VDD(VPWR),
    .Y(_1094_),
    .A(net842),
    .VSS(VGND));
 sg13g2_inv_1 _1744_ (.VDD(VPWR),
    .Y(_1095_),
    .A(net854),
    .VSS(VGND));
 sg13g2_inv_1 _1745_ (.VDD(VPWR),
    .Y(_1096_),
    .A(net844),
    .VSS(VGND));
 sg13g2_inv_1 _1746_ (.VDD(VPWR),
    .Y(_1097_),
    .A(net829),
    .VSS(VGND));
 sg13g2_inv_1 _1747_ (.VDD(VPWR),
    .Y(_1098_),
    .A(net755),
    .VSS(VGND));
 sg13g2_inv_1 _1748_ (.VDD(VPWR),
    .Y(_1099_),
    .A(net711),
    .VSS(VGND));
 sg13g2_inv_1 _1749_ (.VDD(VPWR),
    .Y(_1100_),
    .A(net843),
    .VSS(VGND));
 sg13g2_inv_1 _1750_ (.VDD(VPWR),
    .Y(_1101_),
    .A(net790),
    .VSS(VGND));
 sg13g2_inv_1 _1751_ (.VDD(VPWR),
    .Y(_1102_),
    .A(net400),
    .VSS(VGND));
 sg13g2_inv_1 _1752_ (.VDD(VPWR),
    .Y(_1103_),
    .A(net682),
    .VSS(VGND));
 sg13g2_inv_1 _1753_ (.VDD(VPWR),
    .Y(_1104_),
    .A(net813),
    .VSS(VGND));
 sg13g2_inv_1 _1754_ (.VDD(VPWR),
    .Y(_1105_),
    .A(net394),
    .VSS(VGND));
 sg13g2_inv_1 _1755_ (.VDD(VPWR),
    .Y(_1106_),
    .A(net380),
    .VSS(VGND));
 sg13g2_inv_1 _1756_ (.VDD(VPWR),
    .Y(_1107_),
    .A(net717),
    .VSS(VGND));
 sg13g2_inv_1 _1757_ (.VDD(VPWR),
    .Y(_1108_),
    .A(net438),
    .VSS(VGND));
 sg13g2_inv_1 _1758_ (.VDD(VPWR),
    .Y(_1109_),
    .A(net834),
    .VSS(VGND));
 sg13g2_inv_1 _1759_ (.VDD(VPWR),
    .Y(_1110_),
    .A(net814),
    .VSS(VGND));
 sg13g2_inv_1 _1760_ (.VDD(VPWR),
    .Y(_1111_),
    .A(net430),
    .VSS(VGND));
 sg13g2_inv_1 _1761_ (.VDD(VPWR),
    .Y(_1112_),
    .A(net846),
    .VSS(VGND));
 sg13g2_inv_1 _1762_ (.VDD(VPWR),
    .Y(_1113_),
    .A(net378),
    .VSS(VGND));
 sg13g2_inv_1 _1763_ (.VDD(VPWR),
    .Y(_1114_),
    .A(net863),
    .VSS(VGND));
 sg13g2_inv_1 _1764_ (.VDD(VPWR),
    .Y(_1115_),
    .A(net848),
    .VSS(VGND));
 sg13g2_inv_1 _1765_ (.VDD(VPWR),
    .Y(_1116_),
    .A(net398),
    .VSS(VGND));
 sg13g2_inv_1 _1766_ (.VDD(VPWR),
    .Y(_1117_),
    .A(net706),
    .VSS(VGND));
 sg13g2_inv_1 _1767_ (.VDD(VPWR),
    .Y(_1118_),
    .A(net733),
    .VSS(VGND));
 sg13g2_inv_1 _1768_ (.VDD(VPWR),
    .Y(_1119_),
    .A(net697),
    .VSS(VGND));
 sg13g2_inv_1 _1769_ (.VDD(VPWR),
    .Y(_1120_),
    .A(net850),
    .VSS(VGND));
 sg13g2_inv_1 _1770_ (.VDD(VPWR),
    .Y(_1121_),
    .A(net699),
    .VSS(VGND));
 sg13g2_inv_1 _1771_ (.VDD(VPWR),
    .Y(_1122_),
    .A(net738),
    .VSS(VGND));
 sg13g2_inv_1 _1772_ (.VDD(VPWR),
    .Y(_1123_),
    .A(net810),
    .VSS(VGND));
 sg13g2_inv_1 _1773_ (.VDD(VPWR),
    .Y(_1124_),
    .A(net825),
    .VSS(VGND));
 sg13g2_inv_1 _1774_ (.VDD(VPWR),
    .Y(_1125_),
    .A(net744),
    .VSS(VGND));
 sg13g2_inv_1 _1775_ (.VDD(VPWR),
    .Y(_1126_),
    .A(net780),
    .VSS(VGND));
 sg13g2_inv_1 _1776_ (.VDD(VPWR),
    .Y(_1127_),
    .A(net753),
    .VSS(VGND));
 sg13g2_inv_1 _1777_ (.VDD(VPWR),
    .Y(_1128_),
    .A(net336),
    .VSS(VGND));
 sg13g2_inv_1 _1778_ (.VDD(VPWR),
    .Y(_1129_),
    .A(net350),
    .VSS(VGND));
 sg13g2_inv_1 _1779_ (.VDD(VPWR),
    .Y(_1130_),
    .A(net425),
    .VSS(VGND));
 sg13g2_inv_1 _1780_ (.VDD(VPWR),
    .Y(_1131_),
    .A(net359),
    .VSS(VGND));
 sg13g2_inv_1 _1781_ (.VDD(VPWR),
    .Y(_1132_),
    .A(net714),
    .VSS(VGND));
 sg13g2_inv_1 _1782_ (.VDD(VPWR),
    .Y(_1133_),
    .A(net732),
    .VSS(VGND));
 sg13g2_inv_1 _1783_ (.VDD(VPWR),
    .Y(_1134_),
    .A(net851),
    .VSS(VGND));
 sg13g2_inv_1 _1784_ (.VDD(VPWR),
    .Y(_1135_),
    .A(net338),
    .VSS(VGND));
 sg13g2_inv_1 _1785_ (.VDD(VPWR),
    .Y(_1136_),
    .A(net402),
    .VSS(VGND));
 sg13g2_inv_1 _1786_ (.VDD(VPWR),
    .Y(_1137_),
    .A(net871),
    .VSS(VGND));
 sg13g2_inv_1 _1787_ (.VDD(VPWR),
    .Y(_1138_),
    .A(net794),
    .VSS(VGND));
 sg13g2_inv_1 _1788_ (.VDD(VPWR),
    .Y(_1139_),
    .A(net867),
    .VSS(VGND));
 sg13g2_inv_1 _1789_ (.VDD(VPWR),
    .Y(_1140_),
    .A(net875),
    .VSS(VGND));
 sg13g2_inv_1 _1790_ (.VDD(VPWR),
    .Y(_1141_),
    .A(net703),
    .VSS(VGND));
 sg13g2_inv_1 _1791_ (.VDD(VPWR),
    .Y(_1142_),
    .A(net823),
    .VSS(VGND));
 sg13g2_inv_1 _1792_ (.VDD(VPWR),
    .Y(_1143_),
    .A(net841),
    .VSS(VGND));
 sg13g2_inv_1 _1793_ (.VDD(VPWR),
    .Y(_1144_),
    .A(net771),
    .VSS(VGND));
 sg13g2_inv_1 _1794_ (.VDD(VPWR),
    .Y(_1145_),
    .A(net797),
    .VSS(VGND));
 sg13g2_inv_1 _1795_ (.VDD(VPWR),
    .Y(_1146_),
    .A(net357),
    .VSS(VGND));
 sg13g2_inv_1 _1796_ (.VDD(VPWR),
    .Y(_1147_),
    .A(net361),
    .VSS(VGND));
 sg13g2_inv_1 _1797_ (.VDD(VPWR),
    .Y(_1148_),
    .A(net735),
    .VSS(VGND));
 sg13g2_inv_1 _1798_ (.VDD(VPWR),
    .Y(_1149_),
    .A(net436),
    .VSS(VGND));
 sg13g2_inv_1 _1799_ (.VDD(VPWR),
    .Y(_1150_),
    .A(net806),
    .VSS(VGND));
 sg13g2_inv_1 _1800_ (.VDD(VPWR),
    .Y(_1151_),
    .A(net679),
    .VSS(VGND));
 sg13g2_inv_1 _1801_ (.VDD(VPWR),
    .Y(_1152_),
    .A(net332),
    .VSS(VGND));
 sg13g2_inv_1 _1802_ (.VDD(VPWR),
    .Y(_1153_),
    .A(net781),
    .VSS(VGND));
 sg13g2_inv_1 _1803_ (.VDD(VPWR),
    .Y(_1154_),
    .A(net368),
    .VSS(VGND));
 sg13g2_inv_1 _1804_ (.VDD(VPWR),
    .Y(_1155_),
    .A(net330),
    .VSS(VGND));
 sg13g2_inv_1 _1805_ (.VDD(VPWR),
    .Y(_1156_),
    .A(net747),
    .VSS(VGND));
 sg13g2_inv_1 _1806_ (.VDD(VPWR),
    .Y(_1157_),
    .A(net411),
    .VSS(VGND));
 sg13g2_inv_1 _1807_ (.VDD(VPWR),
    .Y(_1158_),
    .A(net355),
    .VSS(VGND));
 sg13g2_inv_1 _1808_ (.VDD(VPWR),
    .Y(_1159_),
    .A(net351),
    .VSS(VGND));
 sg13g2_inv_1 _1809_ (.VDD(VPWR),
    .Y(_1160_),
    .A(net435),
    .VSS(VGND));
 sg13g2_inv_1 _1810_ (.VDD(VPWR),
    .Y(_1161_),
    .A(net668),
    .VSS(VGND));
 sg13g2_inv_1 _1811_ (.VDD(VPWR),
    .Y(_1162_),
    .A(net428),
    .VSS(VGND));
 sg13g2_inv_1 _1812_ (.VDD(VPWR),
    .Y(_1163_),
    .A(net384),
    .VSS(VGND));
 sg13g2_inv_1 _1813_ (.VDD(VPWR),
    .Y(_1164_),
    .A(net692),
    .VSS(VGND));
 sg13g2_inv_1 _1814_ (.VDD(VPWR),
    .Y(_1165_),
    .A(net831),
    .VSS(VGND));
 sg13g2_inv_1 _1815_ (.VDD(VPWR),
    .Y(_1166_),
    .A(net405),
    .VSS(VGND));
 sg13g2_inv_1 _1816_ (.VDD(VPWR),
    .Y(_1167_),
    .A(net340),
    .VSS(VGND));
 sg13g2_inv_1 _1817_ (.VDD(VPWR),
    .Y(_1168_),
    .A(net773),
    .VSS(VGND));
 sg13g2_inv_1 _1818_ (.VDD(VPWR),
    .Y(_1169_),
    .A(net798),
    .VSS(VGND));
 sg13g2_inv_1 _1819_ (.VDD(VPWR),
    .Y(_1170_),
    .A(net666),
    .VSS(VGND));
 sg13g2_inv_1 _1820_ (.VDD(VPWR),
    .Y(_1171_),
    .A(net382),
    .VSS(VGND));
 sg13g2_inv_1 _1821_ (.VDD(VPWR),
    .Y(_1172_),
    .A(net746),
    .VSS(VGND));
 sg13g2_inv_1 _1822_ (.VDD(VPWR),
    .Y(_1173_),
    .A(net742),
    .VSS(VGND));
 sg13g2_inv_1 _1823_ (.VDD(VPWR),
    .Y(_1174_),
    .A(net362),
    .VSS(VGND));
 sg13g2_inv_1 _1824_ (.VDD(VPWR),
    .Y(_1175_),
    .A(net737),
    .VSS(VGND));
 sg13g2_inv_1 _1825_ (.VDD(VPWR),
    .Y(_1176_),
    .A(net760),
    .VSS(VGND));
 sg13g2_inv_1 _1826_ (.VDD(VPWR),
    .Y(_1177_),
    .A(net839),
    .VSS(VGND));
 sg13g2_inv_1 _1827_ (.VDD(VPWR),
    .Y(_1178_),
    .A(net768),
    .VSS(VGND));
 sg13g2_inv_1 _1828_ (.VDD(VPWR),
    .Y(_1179_),
    .A(net779),
    .VSS(VGND));
 sg13g2_inv_1 _1829_ (.VDD(VPWR),
    .Y(_1180_),
    .A(net673),
    .VSS(VGND));
 sg13g2_inv_1 _1830_ (.VDD(VPWR),
    .Y(_1181_),
    .A(net819),
    .VSS(VGND));
 sg13g2_inv_1 _1831_ (.VDD(VPWR),
    .Y(_1182_),
    .A(net763),
    .VSS(VGND));
 sg13g2_inv_1 _1832_ (.VDD(VPWR),
    .Y(_1183_),
    .A(net386),
    .VSS(VGND));
 sg13g2_inv_1 _1833_ (.VDD(VPWR),
    .Y(_1184_),
    .A(net757),
    .VSS(VGND));
 sg13g2_inv_1 _1834_ (.VDD(VPWR),
    .Y(_1185_),
    .A(net730),
    .VSS(VGND));
 sg13g2_inv_1 _1835_ (.VDD(VPWR),
    .Y(_1186_),
    .A(net828),
    .VSS(VGND));
 sg13g2_inv_1 _1836_ (.VDD(VPWR),
    .Y(_1187_),
    .A(net855),
    .VSS(VGND));
 sg13g2_inv_1 _1837_ (.VDD(VPWR),
    .Y(_1188_),
    .A(net859),
    .VSS(VGND));
 sg13g2_inv_1 _1838_ (.VDD(VPWR),
    .Y(_1189_),
    .A(net775),
    .VSS(VGND));
 sg13g2_inv_1 _1839_ (.VDD(VPWR),
    .Y(_1190_),
    .A(net416),
    .VSS(VGND));
 sg13g2_inv_1 _1840_ (.VDD(VPWR),
    .Y(_1191_),
    .A(net805),
    .VSS(VGND));
 sg13g2_inv_1 _1841_ (.VDD(VPWR),
    .Y(_1192_),
    .A(net388),
    .VSS(VGND));
 sg13g2_inv_1 _1842_ (.VDD(VPWR),
    .Y(_1193_),
    .A(net868),
    .VSS(VGND));
 sg13g2_inv_1 _1843_ (.VDD(VPWR),
    .Y(_1194_),
    .A(net865),
    .VSS(VGND));
 sg13g2_inv_1 _1844_ (.VDD(VPWR),
    .Y(_1195_),
    .A(net860),
    .VSS(VGND));
 sg13g2_inv_1 _1845_ (.VDD(VPWR),
    .Y(_1196_),
    .A(net836),
    .VSS(VGND));
 sg13g2_inv_1 _1846_ (.VDD(VPWR),
    .Y(_1197_),
    .A(net816),
    .VSS(VGND));
 sg13g2_inv_1 _1847_ (.VDD(VPWR),
    .Y(_1198_),
    .A(net708),
    .VSS(VGND));
 sg13g2_inv_1 _1848_ (.VDD(VPWR),
    .Y(_1199_),
    .A(net421),
    .VSS(VGND));
 sg13g2_inv_1 _1849_ (.VDD(VPWR),
    .Y(_1200_),
    .A(net739),
    .VSS(VGND));
 sg13g2_inv_1 _1850_ (.VDD(VPWR),
    .Y(_1201_),
    .A(net821),
    .VSS(VGND));
 sg13g2_inv_1 _1851_ (.VDD(VPWR),
    .Y(_1202_),
    .A(net801),
    .VSS(VGND));
 sg13g2_inv_1 _1852_ (.VDD(VPWR),
    .Y(_1203_),
    .A(net342),
    .VSS(VGND));
 sg13g2_inv_1 _1853_ (.VDD(VPWR),
    .Y(_1204_),
    .A(net684),
    .VSS(VGND));
 sg13g2_inv_1 _1854_ (.VDD(VPWR),
    .Y(_1205_),
    .A(net442),
    .VSS(VGND));
 sg13g2_inv_1 _1855_ (.VDD(VPWR),
    .Y(_1206_),
    .A(net423),
    .VSS(VGND));
 sg13g2_inv_1 _1856_ (.VDD(VPWR),
    .Y(_1207_),
    .A(net770),
    .VSS(VGND));
 sg13g2_inv_1 _1857_ (.VDD(VPWR),
    .Y(_1208_),
    .A(net370),
    .VSS(VGND));
 sg13g2_inv_1 _1858_ (.VDD(VPWR),
    .Y(_1209_),
    .A(net789),
    .VSS(VGND));
 sg13g2_inv_1 _1859_ (.VDD(VPWR),
    .Y(_1210_),
    .A(net784),
    .VSS(VGND));
 sg13g2_inv_1 _1860_ (.VDD(VPWR),
    .Y(_1211_),
    .A(net796),
    .VSS(VGND));
 sg13g2_inv_1 _1861_ (.VDD(VPWR),
    .Y(_1212_),
    .A(net724),
    .VSS(VGND));
 sg13g2_inv_1 _1862_ (.VDD(VPWR),
    .Y(_1213_),
    .A(net778),
    .VSS(VGND));
 sg13g2_inv_1 _1863_ (.VDD(VPWR),
    .Y(_1214_),
    .A(net677),
    .VSS(VGND));
 sg13g2_inv_1 _1864_ (.VDD(VPWR),
    .Y(_1215_),
    .A(net705),
    .VSS(VGND));
 sg13g2_nor2b_1 _1865_ (.A(net534),
    .B_N(net535),
    .Y(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1866_ (.A(\controller.inst_mem.addr[2] ),
    .B(_1216_),
    .X(_1217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _1867_ (.B(net536),
    .C(net532),
    .Y(_1218_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net533));
 sg13g2_nand2_1 _1868_ (.Y(_1219_),
    .A(\controller.inst_mem.mem_data[159] ),
    .B(net510),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1869_ (.A(_1068_),
    .B(_1216_),
    .X(_1220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _1870_ (.Y(_1221_),
    .B(net533),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net535));
 sg13g2_nor2_1 _1871_ (.A(_1068_),
    .B(_1221_),
    .Y(_1222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _1872_ (.B(net534),
    .C(net531),
    .Y(_1223_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net535));
 sg13g2_a22oi_1 _1873_ (.Y(_1224_),
    .B1(net502),
    .B2(\controller.inst_mem.mem_data[183] ),
    .A2(net506),
    .A1(\controller.inst_mem.mem_data[63] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1874_ (.Y(_1225_),
    .A(net534),
    .B(net535),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1875_ (.A(net531),
    .B(_1225_),
    .Y(_1226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1876_ (.A(net531),
    .B(_1221_),
    .Y(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1877_ (.Y(_1228_),
    .B1(net494),
    .B2(\controller.inst_mem.mem_data[87] ),
    .A2(net498),
    .A1(\controller.inst_mem.mem_data[111] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _1878_ (.X(_1229_),
    .A(net532),
    .B(net533),
    .C(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1879_ (.A(net533),
    .B(net536),
    .Y(_1230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _1880_ (.A(net532),
    .B(net533),
    .C(net536),
    .Y(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1881_ (.Y(_1232_),
    .A(_1068_),
    .B(net520),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1882_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[135] ),
    .C1(net514),
    .B1(net519),
    .A1(\controller.inst_mem.extended_word[7] ),
    .Y(_1233_),
    .A2(net523));
 sg13g2_nand4_1 _1883_ (.B(_1224_),
    .C(_1228_),
    .A(_1219_),
    .Y(_1234_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1233_));
 sg13g2_o21ai_1 _1884_ (.B1(_1234_),
    .VDD(VPWR),
    .Y(_1235_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[39] ),
    .A2(net493));
 sg13g2_inv_1 _1885_ (.VDD(VPWR),
    .Y(_1236_),
    .A(_1235_),
    .VSS(VGND));
 sg13g2_nand2_1 _1886_ (.Y(_1237_),
    .A(\controller.inst_mem.mem_data[64] ),
    .B(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1887_ (.Y(_1238_),
    .B1(net494),
    .B2(\controller.inst_mem.mem_data[88] ),
    .A2(net502),
    .A1(\controller.inst_mem.mem_data[184] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1888_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[136] ),
    .C1(net514),
    .B1(net519),
    .A1(\controller.inst_mem.mem_data[112] ),
    .Y(_1239_),
    .A2(net498));
 sg13g2_nand2_1 _1889_ (.Y(_1240_),
    .A(_1237_),
    .B(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1890_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.extended_word[8] ),
    .C1(_1240_),
    .B1(net523),
    .A1(\controller.inst_mem.mem_data[160] ),
    .Y(_1241_),
    .A2(net510));
 sg13g2_a22oi_1 _1891_ (.Y(_1242_),
    .B1(_1238_),
    .B2(_1241_),
    .A2(net514),
    .A1(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1892_ (.Y(_1243_),
    .B1(net523),
    .B2(\controller.inst_mem.extended_word[5] ),
    .A2(net494),
    .A1(\controller.inst_mem.mem_data[85] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1893_ (.Y(_1244_),
    .B1(net502),
    .B2(\controller.inst_mem.mem_data[181] ),
    .A2(net510),
    .A1(\controller.inst_mem.mem_data[157] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1894_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[133] ),
    .C1(net514),
    .B1(net519),
    .A1(\controller.inst_mem.mem_data[109] ),
    .Y(_1245_),
    .A2(net498));
 sg13g2_nand3_1 _1895_ (.B(_1244_),
    .C(_1245_),
    .A(_1243_),
    .Y(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1896_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[61] ),
    .A2(net506),
    .Y(_1247_),
    .B1(_1246_));
 sg13g2_a21oi_1 _1897_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1023_),
    .A2(net514),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_inv_1 _1898_ (.VDD(VPWR),
    .Y(_1249_),
    .A(_1248_),
    .VSS(VGND));
 sg13g2_a221oi_1 _1899_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[134] ),
    .C1(net514),
    .B1(net519),
    .A1(\controller.inst_mem.mem_data[86] ),
    .Y(_1250_),
    .A2(net494));
 sg13g2_a22oi_1 _1900_ (.Y(_1251_),
    .B1(net502),
    .B2(\controller.inst_mem.mem_data[182] ),
    .A2(net510),
    .A1(\controller.inst_mem.mem_data[158] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1901_ (.Y(_1252_),
    .B1(net498),
    .B2(\controller.inst_mem.mem_data[110] ),
    .A2(net506),
    .A1(\controller.inst_mem.mem_data[62] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1902_ (.B(_1251_),
    .C(_1252_),
    .A(_1250_),
    .Y(_1253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1903_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.extended_word[6] ),
    .A2(net523),
    .Y(_1254_),
    .B1(_1253_));
 sg13g2_a21o_1 _1904_ (.A2(net514),
    .A1(_1022_),
    .B1(_1254_),
    .X(_1255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1905_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1256_),
    .B(_1255_),
    .A(_1249_));
 sg13g2_or2_1 _1906_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1257_),
    .B(_1256_),
    .A(_1242_));
 sg13g2_nor2_2 _1907_ (.A(_1236_),
    .B(_1257_),
    .Y(_1258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1248_),
    .A2(_1255_),
    .Y(_1259_),
    .B1(_1258_));
 sg13g2_nor2_2 _1909_ (.A(_1235_),
    .B(_1257_),
    .Y(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1910_ (.A(_1235_),
    .B_N(_1242_),
    .Y(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1911_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.output_controller.keep[0] ),
    .A2(_1261_),
    .Y(_1262_),
    .B1(_1249_));
 sg13g2_nor2_1 _1912_ (.A(_1255_),
    .B(_1262_),
    .Y(_1263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1913_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net965),
    .A2(_1260_),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_o21ai_1 _1914_ (.B1(_1264_),
    .VDD(VPWR),
    .Y(net15),
    .VSS(VGND),
    .A1(_1067_),
    .A2(_1259_));
 sg13g2_a22oi_1 _1915_ (.Y(_1265_),
    .B1(_1261_),
    .B2(net940),
    .A2(_1256_),
    .A1(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1916_ (.Y(_1266_),
    .B1(_1260_),
    .B2(\controller.alu_buffer.buffer[17] ),
    .A2(_1258_),
    .A1(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1917_ (.Y(net16),
    .A(_1265_),
    .B(_1266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1918_ (.Y(_1267_),
    .B1(_1261_),
    .B2(net917),
    .A2(_1256_),
    .A1(_1242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1919_ (.Y(_1268_),
    .B1(_1260_),
    .B2(\controller.alu_buffer.buffer[18] ),
    .A2(_1258_),
    .A1(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1920_ (.Y(net17),
    .A(_1267_),
    .B(_1268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1921_ (.A(net911),
    .B(\controller.counter2.counter_1[1] ),
    .C(net892),
    .Y(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _1922_ (.A(\controller.counter2.counter_1[3] ),
    .B(\controller.counter2.counter_1[2] ),
    .C(\controller.counter2.counter_1[1] ),
    .D(\controller.counter2.counter_1[0] ),
    .X(_1270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1923_ (.A(net910),
    .B(net903),
    .C(_1270_),
    .X(_1271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _1924_ (.A(\controller.counter2.counter_1[6] ),
    .B(\controller.counter2.counter_1[5] ),
    .C(\controller.counter2.counter_1[4] ),
    .D(_1270_),
    .X(_1272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1925_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1273_),
    .B(_1272_),
    .A(net932));
 sg13g2_nor4_2 _1926_ (.A(net901),
    .B(\controller.counter2.counter_1[8] ),
    .C(\controller.counter2.counter_1[7] ),
    .Y(_1274_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1272_));
 sg13g2_nand2b_1 _1927_ (.Y(_1275_),
    .B(_1274_),
    .A_N(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1928_ (.A(net883),
    .B(\controller.counter2.counter_1[10] ),
    .Y(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1929_ (.Y(_1277_),
    .A(_1274_),
    .B(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _1930_ (.A(\controller.counter2.counter_1[15] ),
    .B(\controller.counter2.counter_1[14] ),
    .C(\controller.counter2.counter_1[13] ),
    .D(\controller.counter2.counter_1[12] ),
    .Y(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _1931_ (.A(_1277_),
    .B_N(_1278_),
    .Y(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1932_ (.B(_1276_),
    .C(_1278_),
    .A(_1274_),
    .Y(_1280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1933_ (.Y(_1281_),
    .A(\controller.alu_buffer.buffer[19] ),
    .B(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1934_ (.Y(_1282_),
    .B1(_1279_),
    .B2(_1257_),
    .A2(_1258_),
    .A1(\controller.alu_buffer.buffer[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1935_ (.Y(net18),
    .A(_1281_),
    .B(_1282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _1936_ (.A(\controller.alu_buffer.buffer[3] ),
    .B(net529),
    .C(net530),
    .Y(_1283_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net971));
 sg13g2_nor2_1 _1937_ (.A(\controller.alu_buffer.buffer[5] ),
    .B(net528),
    .Y(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1938_ (.Y(_1285_),
    .A(_1283_),
    .B(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1939_ (.A(\controller.alu_buffer.buffer[7] ),
    .B(net527),
    .Y(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1940_ (.B(_1284_),
    .C(_1286_),
    .A(_1283_),
    .Y(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1941_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1288_),
    .B(_1287_),
    .A(\controller.alu_buffer.buffer[8] ));
 sg13g2_nor3_1 _1942_ (.A(\controller.alu_buffer.buffer[10] ),
    .B(\controller.alu_buffer.buffer[9] ),
    .C(\controller.alu_buffer.buffer[8] ),
    .Y(_1289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1943_ (.B(_1284_),
    .C(_1286_),
    .A(_1283_),
    .Y(_1290_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1289_));
 sg13g2_or2_1 _1944_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1291_),
    .B(_1290_),
    .A(\controller.alu_buffer.buffer[11] ));
 sg13g2_nor3_1 _1945_ (.A(\controller.alu_buffer.buffer[14] ),
    .B(\controller.alu_buffer.buffer[13] ),
    .C(\controller.alu_buffer.buffer[12] ),
    .Y(_1292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1946_ (.Y(_1293_),
    .A(_1064_),
    .B(_1292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1947_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1294_),
    .B(_1293_),
    .A(_1291_));
 sg13g2_or4_1 _1948_ (.A(\controller.alu_buffer.buffer[19] ),
    .B(\controller.alu_buffer.buffer[18] ),
    .C(\controller.alu_buffer.buffer[17] ),
    .D(\controller.alu_buffer.buffer[16] ),
    .X(_1295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _1949_ (.A(\controller.alu_buffer.buffer[11] ),
    .B(_1290_),
    .C(_1293_),
    .Y(_1296_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1295_));
 sg13g2_nand2b_1 _1950_ (.Y(_1297_),
    .B(_1296_),
    .A_N(\controller.alu_buffer.buffer[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1951_ (.A(\controller.alu_buffer.buffer[23] ),
    .B(\controller.alu_buffer.buffer[22] ),
    .C(\controller.alu_buffer.buffer[21] ),
    .Y(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1952_ (.A(_1297_),
    .B_N(_1298_),
    .Y(_1299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _1953_ (.B(_1296_),
    .C(_1298_),
    .Y(_1300_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\controller.alu_buffer.buffer[20] ));
 sg13g2_nand2_1 _1954_ (.Y(_1301_),
    .A(\controller.alu_buffer.buffer[20] ),
    .B(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1955_ (.Y(_1302_),
    .B1(_1299_),
    .B2(_1257_),
    .A2(_1258_),
    .A1(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1956_ (.Y(net19),
    .A(_1301_),
    .B(_1302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1957_ (.Y(_1303_),
    .A(\controller.alu_buffer.buffer[21] ),
    .B(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1958_ (.Y(_1304_),
    .B1(_1258_),
    .B2(\controller.alu_buffer.buffer[5] ),
    .A2(_1257_),
    .A1(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1959_ (.Y(net20),
    .A(_1303_),
    .B(_1304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1960_ (.Y(_1305_),
    .A(\controller.alu_buffer.buffer[22] ),
    .B(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1961_ (.Y(_1306_),
    .B1(_1258_),
    .B2(net527),
    .A2(_1257_),
    .A1(net533),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1962_ (.Y(net21),
    .A(_1305_),
    .B(_1306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1963_ (.Y(_1307_),
    .A(\controller.alu_buffer.buffer[23] ),
    .B(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1964_ (.Y(_1308_),
    .B1(_1258_),
    .B2(\controller.alu_buffer.buffer[7] ),
    .A2(_1257_),
    .A1(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1965_ (.Y(net22),
    .A(_1307_),
    .B(_1308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1966_ (.A(net6),
    .B(net5),
    .X(_1309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1967_ (.B1(net643),
    .VDD(VPWR),
    .Y(_1310_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[81] ),
    .A2(net586));
 sg13g2_a21oi_1 _1968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0980_),
    .A2(net586),
    .Y(_0000_),
    .B1(_1310_));
 sg13g2_o21ai_1 _1969_ (.B1(net643),
    .VDD(VPWR),
    .Y(_1311_),
    .VSS(VGND),
    .A1(net677),
    .A2(net586));
 sg13g2_a21oi_1 _1970_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1215_),
    .A2(net586),
    .Y(_0001_),
    .B1(_1311_));
 sg13g2_o21ai_1 _1971_ (.B1(net642),
    .VDD(VPWR),
    .Y(_1312_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[83] ),
    .A2(net581));
 sg13g2_a21oi_1 _1972_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1214_),
    .A2(net581),
    .Y(_0002_),
    .B1(_1312_));
 sg13g2_o21ai_1 _1973_ (.B1(net630),
    .VDD(VPWR),
    .Y(_1313_),
    .VSS(VGND),
    .A1(net724),
    .A2(net559));
 sg13g2_a21oi_1 _1974_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1213_),
    .A2(net559),
    .Y(_0003_),
    .B1(_1313_));
 sg13g2_o21ai_1 _1975_ (.B1(net628),
    .VDD(VPWR),
    .Y(_1314_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[85] ),
    .A2(net555));
 sg13g2_a21oi_1 _1976_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1212_),
    .A2(net555),
    .Y(_0004_),
    .B1(_1314_));
 sg13g2_o21ai_1 _1977_ (.B1(net628),
    .VDD(VPWR),
    .Y(_1315_),
    .VSS(VGND),
    .A1(net784),
    .A2(net550));
 sg13g2_a21oi_1 _1978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1211_),
    .A2(net557),
    .Y(_0005_),
    .B1(_1315_));
 sg13g2_o21ai_1 _1979_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1316_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[87] ),
    .A2(net548));
 sg13g2_a21oi_1 _1980_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1210_),
    .A2(net548),
    .Y(_0006_),
    .B1(_1316_));
 sg13g2_o21ai_1 _1981_ (.B1(net626),
    .VDD(VPWR),
    .Y(_1317_),
    .VSS(VGND),
    .A1(net370),
    .A2(net551));
 sg13g2_a21oi_1 _1982_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1209_),
    .A2(net546),
    .Y(_0007_),
    .B1(_1317_));
 sg13g2_o21ai_1 _1983_ (.B1(net629),
    .VDD(VPWR),
    .Y(_1318_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[89] ),
    .A2(net552));
 sg13g2_a21oi_1 _1984_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1208_),
    .A2(net552),
    .Y(_0008_),
    .B1(_1318_));
 sg13g2_o21ai_1 _1985_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1319_),
    .VSS(VGND),
    .A1(net423),
    .A2(net562));
 sg13g2_a21oi_1 _1986_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1207_),
    .A2(net564),
    .Y(_0009_),
    .B1(_1319_));
 sg13g2_o21ai_1 _1987_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1320_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[91] ),
    .A2(net566));
 sg13g2_a21oi_1 _1988_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1206_),
    .A2(net566),
    .Y(_0010_),
    .B1(_1320_));
 sg13g2_o21ai_1 _1989_ (.B1(net633),
    .VDD(VPWR),
    .Y(_1321_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[92] ),
    .A2(net567));
 sg13g2_a21oi_1 _1990_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1205_),
    .A2(net567),
    .Y(_0011_),
    .B1(_1321_));
 sg13g2_o21ai_1 _1991_ (.B1(net655),
    .VDD(VPWR),
    .Y(_1322_),
    .VSS(VGND),
    .A1(net342),
    .A2(net607));
 sg13g2_a21oi_1 _1992_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1204_),
    .A2(net572),
    .Y(_0012_),
    .B1(_1322_));
 sg13g2_o21ai_1 _1993_ (.B1(net655),
    .VDD(VPWR),
    .Y(_1323_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[94] ),
    .A2(net607));
 sg13g2_a21oi_1 _1994_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1203_),
    .A2(net607),
    .Y(_0013_),
    .B1(_1323_));
 sg13g2_o21ai_1 _1995_ (.B1(net656),
    .VDD(VPWR),
    .Y(_1324_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[95] ),
    .A2(net610));
 sg13g2_a21oi_1 _1996_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1202_),
    .A2(net609),
    .Y(_0014_),
    .B1(_1324_));
 sg13g2_o21ai_1 _1997_ (.B1(net660),
    .VDD(VPWR),
    .Y(_1325_),
    .VSS(VGND),
    .A1(net739),
    .A2(net617));
 sg13g2_a21oi_1 _1998_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1201_),
    .A2(net617),
    .Y(_0015_),
    .B1(_1325_));
 sg13g2_o21ai_1 _1999_ (.B1(net662),
    .VDD(VPWR),
    .Y(_1326_),
    .VSS(VGND),
    .A1(net421),
    .A2(net618));
 sg13g2_a21oi_1 _2000_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1200_),
    .A2(net618),
    .Y(_0016_),
    .B1(_1326_));
 sg13g2_o21ai_1 _2001_ (.B1(net661),
    .VDD(VPWR),
    .Y(_1327_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[98] ),
    .A2(net619));
 sg13g2_a21oi_1 _2002_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1199_),
    .A2(net619),
    .Y(_0017_),
    .B1(_1327_));
 sg13g2_o21ai_1 _2003_ (.B1(net651),
    .VDD(VPWR),
    .Y(_1328_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[99] ),
    .A2(net601));
 sg13g2_a21oi_1 _2004_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1198_),
    .A2(net620),
    .Y(_0018_),
    .B1(_1328_));
 sg13g2_o21ai_1 _2005_ (.B1(net651),
    .VDD(VPWR),
    .Y(_1329_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[100] ),
    .A2(net601));
 sg13g2_a21oi_1 _2006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1197_),
    .A2(net601),
    .Y(_0019_),
    .B1(_1329_));
 sg13g2_o21ai_1 _2007_ (.B1(net652),
    .VDD(VPWR),
    .Y(_1330_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[101] ),
    .A2(net600));
 sg13g2_a21oi_1 _2008_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1196_),
    .A2(net600),
    .Y(_0020_),
    .B1(_1330_));
 sg13g2_o21ai_1 _2009_ (.B1(net649),
    .VDD(VPWR),
    .Y(_1331_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[102] ),
    .A2(net595));
 sg13g2_a21oi_1 _2010_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1195_),
    .A2(net595),
    .Y(_0021_),
    .B1(_1331_));
 sg13g2_o21ai_1 _2011_ (.B1(net649),
    .VDD(VPWR),
    .Y(_1332_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[103] ),
    .A2(net595));
 sg13g2_a21oi_1 _2012_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1194_),
    .A2(net595),
    .Y(_0022_),
    .B1(_1332_));
 sg13g2_o21ai_1 _2013_ (.B1(net649),
    .VDD(VPWR),
    .Y(_1333_),
    .VSS(VGND),
    .A1(net388),
    .A2(net597));
 sg13g2_a21oi_1 _2014_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1193_),
    .A2(net597),
    .Y(_0023_),
    .B1(_1333_));
 sg13g2_o21ai_1 _2015_ (.B1(net648),
    .VDD(VPWR),
    .Y(_1334_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[105] ),
    .A2(net592));
 sg13g2_a21oi_1 _2016_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1192_),
    .A2(net592),
    .Y(_0024_),
    .B1(_1334_));
 sg13g2_o21ai_1 _2017_ (.B1(net643),
    .VDD(VPWR),
    .Y(_1335_),
    .VSS(VGND),
    .A1(net416),
    .A2(net585));
 sg13g2_a21oi_1 _2018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1191_),
    .A2(net585),
    .Y(_0025_),
    .B1(_1335_));
 sg13g2_o21ai_1 _2019_ (.B1(net642),
    .VDD(VPWR),
    .Y(_1336_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[107] ),
    .A2(net581));
 sg13g2_a21oi_1 _2020_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1190_),
    .A2(net581),
    .Y(_0026_),
    .B1(_1336_));
 sg13g2_o21ai_1 _2021_ (.B1(net630),
    .VDD(VPWR),
    .Y(_1337_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[108] ),
    .A2(net559));
 sg13g2_a21oi_1 _2022_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1189_),
    .A2(net559),
    .Y(_0027_),
    .B1(_1337_));
 sg13g2_o21ai_1 _2023_ (.B1(net628),
    .VDD(VPWR),
    .Y(_1338_),
    .VSS(VGND),
    .A1(net855),
    .A2(net555));
 sg13g2_a21oi_1 _2024_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1188_),
    .A2(net555),
    .Y(_0028_),
    .B1(_1338_));
 sg13g2_o21ai_1 _2025_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1339_),
    .VSS(VGND),
    .A1(net828),
    .A2(net550));
 sg13g2_a21oi_1 _2026_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1187_),
    .A2(net550),
    .Y(_0029_),
    .B1(_1339_));
 sg13g2_o21ai_1 _2027_ (.B1(net625),
    .VDD(VPWR),
    .Y(_0289_),
    .VSS(VGND),
    .A1(net730),
    .A2(net549));
 sg13g2_a21oi_1 _2028_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1186_),
    .A2(net548),
    .Y(_0030_),
    .B1(_0289_));
 sg13g2_o21ai_1 _2029_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0290_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[112] ),
    .A2(net552));
 sg13g2_a21oi_1 _2030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1185_),
    .A2(net550),
    .Y(_0031_),
    .B1(_0290_));
 sg13g2_o21ai_1 _2031_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0291_),
    .VSS(VGND),
    .A1(net386),
    .A2(net558));
 sg13g2_a21oi_1 _2032_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1184_),
    .A2(net558),
    .Y(_0032_),
    .B1(_0291_));
 sg13g2_o21ai_1 _2033_ (.B1(net633),
    .VDD(VPWR),
    .Y(_0292_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[114] ),
    .A2(net566));
 sg13g2_a21oi_1 _2034_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1183_),
    .A2(net566),
    .Y(_0033_),
    .B1(_0292_));
 sg13g2_o21ai_1 _2035_ (.B1(net633),
    .VDD(VPWR),
    .Y(_0293_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[115] ),
    .A2(net566));
 sg13g2_a21oi_1 _2036_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1182_),
    .A2(net566),
    .Y(_0034_),
    .B1(_0293_));
 sg13g2_o21ai_1 _2037_ (.B1(net634),
    .VDD(VPWR),
    .Y(_0294_),
    .VSS(VGND),
    .A1(net673),
    .A2(net565));
 sg13g2_a21oi_1 _2038_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1181_),
    .A2(net565),
    .Y(_0035_),
    .B1(_0294_));
 sg13g2_o21ai_1 _2039_ (.B1(net655),
    .VDD(VPWR),
    .Y(_0295_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[117] ),
    .A2(net573));
 sg13g2_a21oi_1 _2040_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1180_),
    .A2(net573),
    .Y(_0036_),
    .B1(_0295_));
 sg13g2_o21ai_1 _2041_ (.B1(net655),
    .VDD(VPWR),
    .Y(_0296_),
    .VSS(VGND),
    .A1(net768),
    .A2(net606));
 sg13g2_a21oi_1 _2042_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1179_),
    .A2(net606),
    .Y(_0037_),
    .B1(_0296_));
 sg13g2_o21ai_1 _2043_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0297_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[119] ),
    .A2(net609));
 sg13g2_a21oi_1 _2044_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1178_),
    .A2(net609),
    .Y(_0038_),
    .B1(_0297_));
 sg13g2_o21ai_1 _2045_ (.B1(net662),
    .VDD(VPWR),
    .Y(_0298_),
    .VSS(VGND),
    .A1(net760),
    .A2(net617));
 sg13g2_a21oi_1 _2046_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1177_),
    .A2(net617),
    .Y(_0039_),
    .B1(_0298_));
 sg13g2_o21ai_1 _2047_ (.B1(net662),
    .VDD(VPWR),
    .Y(_0299_),
    .VSS(VGND),
    .A1(net737),
    .A2(net621));
 sg13g2_a21oi_1 _2048_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1176_),
    .A2(net618),
    .Y(_0040_),
    .B1(_0299_));
 sg13g2_o21ai_1 _2049_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0300_),
    .VSS(VGND),
    .A1(net362),
    .A2(net621));
 sg13g2_a21oi_1 _2050_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1175_),
    .A2(net621),
    .Y(_0041_),
    .B1(_0300_));
 sg13g2_o21ai_1 _2051_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0301_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[123] ),
    .A2(net620));
 sg13g2_a21oi_1 _2052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1174_),
    .A2(net620),
    .Y(_0042_),
    .B1(_0301_));
 sg13g2_o21ai_1 _2053_ (.B1(net651),
    .VDD(VPWR),
    .Y(_0302_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[124] ),
    .A2(net602));
 sg13g2_a21oi_1 _2054_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1173_),
    .A2(net602),
    .Y(_0043_),
    .B1(_0302_));
 sg13g2_o21ai_1 _2055_ (.B1(net652),
    .VDD(VPWR),
    .Y(_0303_),
    .VSS(VGND),
    .A1(net382),
    .A2(net599));
 sg13g2_a21oi_1 _2056_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1172_),
    .A2(net599),
    .Y(_0044_),
    .B1(_0303_));
 sg13g2_o21ai_1 _2057_ (.B1(net649),
    .VDD(VPWR),
    .Y(_0304_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[126] ),
    .A2(net596));
 sg13g2_a21oi_1 _2058_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1171_),
    .A2(net596),
    .Y(_0045_),
    .B1(_0304_));
 sg13g2_o21ai_1 _2059_ (.B1(net650),
    .VDD(VPWR),
    .Y(_0305_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[127] ),
    .A2(net596));
 sg13g2_a21oi_1 _2060_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1170_),
    .A2(net596),
    .Y(_0046_),
    .B1(_0305_));
 sg13g2_o21ai_1 _2061_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0306_),
    .VSS(VGND),
    .A1(net773),
    .A2(net592));
 sg13g2_a21oi_1 _2062_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1169_),
    .A2(net592),
    .Y(_0047_),
    .B1(_0306_));
 sg13g2_o21ai_1 _2063_ (.B1(net643),
    .VDD(VPWR),
    .Y(_0307_),
    .VSS(VGND),
    .A1(net340),
    .A2(net587));
 sg13g2_a21oi_1 _2064_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1168_),
    .A2(net586),
    .Y(_0048_),
    .B1(_0307_));
 sg13g2_o21ai_1 _2065_ (.B1(net643),
    .VDD(VPWR),
    .Y(_0308_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[130] ),
    .A2(net585));
 sg13g2_a21oi_1 _2066_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1167_),
    .A2(net585),
    .Y(_0049_),
    .B1(_0308_));
 sg13g2_o21ai_1 _2067_ (.B1(net642),
    .VDD(VPWR),
    .Y(_0309_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[131] ),
    .A2(net581));
 sg13g2_a21oi_1 _2068_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1166_),
    .A2(net584),
    .Y(_0050_),
    .B1(_0309_));
 sg13g2_o21ai_1 _2069_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0310_),
    .VSS(VGND),
    .A1(net692),
    .A2(net560));
 sg13g2_a21oi_1 _2070_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1165_),
    .A2(net560),
    .Y(_0051_),
    .B1(_0310_));
 sg13g2_o21ai_1 _2071_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0311_),
    .VSS(VGND),
    .A1(net384),
    .A2(net556));
 sg13g2_a21oi_1 _2072_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1164_),
    .A2(net556),
    .Y(_0052_),
    .B1(_0311_));
 sg13g2_o21ai_1 _2073_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0312_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[134] ),
    .A2(net557));
 sg13g2_a21oi_1 _2074_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1163_),
    .A2(net557),
    .Y(_0053_),
    .B1(_0312_));
 sg13g2_o21ai_1 _2075_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0313_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[135] ),
    .A2(net550));
 sg13g2_a21oi_1 _2076_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1162_),
    .A2(net550),
    .Y(_0054_),
    .B1(_0313_));
 sg13g2_o21ai_1 _2077_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0314_),
    .VSS(VGND),
    .A1(net435),
    .A2(net552));
 sg13g2_a21oi_1 _2078_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1161_),
    .A2(net552),
    .Y(_0055_),
    .B1(_0314_));
 sg13g2_o21ai_1 _2079_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0315_),
    .VSS(VGND),
    .A1(net351),
    .A2(net558));
 sg13g2_a21oi_1 _2080_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1160_),
    .A2(net558),
    .Y(_0056_),
    .B1(_0315_));
 sg13g2_o21ai_1 _2081_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0316_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[138] ),
    .A2(net562));
 sg13g2_a21oi_1 _2082_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1159_),
    .A2(net562),
    .Y(_0057_),
    .B1(_0316_));
 sg13g2_o21ai_1 _2083_ (.B1(net633),
    .VDD(VPWR),
    .Y(_0317_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[139] ),
    .A2(net566));
 sg13g2_a21oi_1 _2084_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1158_),
    .A2(net566),
    .Y(_0058_),
    .B1(_0317_));
 sg13g2_o21ai_1 _2085_ (.B1(net633),
    .VDD(VPWR),
    .Y(_0318_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[140] ),
    .A2(net565));
 sg13g2_a21oi_1 _2086_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1157_),
    .A2(net565),
    .Y(_0059_),
    .B1(_0318_));
 sg13g2_o21ai_1 _2087_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0319_),
    .VSS(VGND),
    .A1(net330),
    .A2(net590));
 sg13g2_a21oi_1 _2088_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1156_),
    .A2(net590),
    .Y(_0060_),
    .B1(_0319_));
 sg13g2_o21ai_1 _2089_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0320_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[142] ),
    .A2(net590));
 sg13g2_a21oi_1 _2090_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1155_),
    .A2(net590),
    .Y(_0061_),
    .B1(_0320_));
 sg13g2_o21ai_1 _2091_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0321_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[143] ),
    .A2(net588));
 sg13g2_a21oi_1 _2092_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1154_),
    .A2(net588),
    .Y(_0062_),
    .B1(_0321_));
 sg13g2_o21ai_1 _2093_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0322_),
    .VSS(VGND),
    .A1(net332),
    .A2(net616));
 sg13g2_a21oi_1 _2094_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1153_),
    .A2(net608),
    .Y(_0063_),
    .B1(_0322_));
 sg13g2_o21ai_1 _2095_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0323_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[145] ),
    .A2(net615));
 sg13g2_a21oi_1 _2096_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1152_),
    .A2(net615),
    .Y(_0064_),
    .B1(_0323_));
 sg13g2_o21ai_1 _2097_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0324_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[146] ),
    .A2(net615));
 sg13g2_a21oi_1 _2098_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1151_),
    .A2(net615),
    .Y(_0065_),
    .B1(_0324_));
 sg13g2_o21ai_1 _2099_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0325_),
    .VSS(VGND),
    .A1(net436),
    .A2(net598));
 sg13g2_a21oi_1 _2100_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1150_),
    .A2(net604),
    .Y(_0066_),
    .B1(_0325_));
 sg13g2_o21ai_1 _2101_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0326_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[148] ),
    .A2(net598));
 sg13g2_a21oi_1 _2102_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1149_),
    .A2(net604),
    .Y(_0067_),
    .B1(_0326_));
 sg13g2_o21ai_1 _2103_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0327_),
    .VSS(VGND),
    .A1(net361),
    .A2(net598));
 sg13g2_a21oi_1 _2104_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1148_),
    .A2(net598),
    .Y(_0068_),
    .B1(_0327_));
 sg13g2_o21ai_1 _2105_ (.B1(net650),
    .VDD(VPWR),
    .Y(_0328_),
    .VSS(VGND),
    .A1(net357),
    .A2(net593));
 sg13g2_a21oi_1 _2106_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1147_),
    .A2(net593),
    .Y(_0069_),
    .B1(_0328_));
 sg13g2_o21ai_1 _2107_ (.B1(net650),
    .VDD(VPWR),
    .Y(_0329_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[151] ),
    .A2(net593));
 sg13g2_a21oi_1 _2108_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1146_),
    .A2(net594),
    .Y(_0070_),
    .B1(_0329_));
 sg13g2_o21ai_1 _2109_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0330_),
    .VSS(VGND),
    .A1(net771),
    .A2(net592));
 sg13g2_a21oi_1 _2110_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1145_),
    .A2(net592),
    .Y(_0071_),
    .B1(_0330_));
 sg13g2_o21ai_1 _2111_ (.B1(net643),
    .VDD(VPWR),
    .Y(_0331_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[153] ),
    .A2(net586));
 sg13g2_a21oi_1 _2112_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1144_),
    .A2(net586),
    .Y(_0072_),
    .B1(_0331_));
 sg13g2_o21ai_1 _2113_ (.B1(net643),
    .VDD(VPWR),
    .Y(_0332_),
    .VSS(VGND),
    .A1(net823),
    .A2(net585));
 sg13g2_a21oi_1 _2114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1143_),
    .A2(net585),
    .Y(_0073_),
    .B1(_0332_));
 sg13g2_o21ai_1 _2115_ (.B1(net642),
    .VDD(VPWR),
    .Y(_0333_),
    .VSS(VGND),
    .A1(net703),
    .A2(net581));
 sg13g2_a21oi_1 _2116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1142_),
    .A2(net581),
    .Y(_0074_),
    .B1(_0333_));
 sg13g2_o21ai_1 _2117_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0334_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[156] ),
    .A2(net559));
 sg13g2_a21oi_1 _2118_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1141_),
    .A2(net559),
    .Y(_0075_),
    .B1(_0334_));
 sg13g2_o21ai_1 _2119_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0335_),
    .VSS(VGND),
    .A1(net867),
    .A2(net555));
 sg13g2_a21oi_1 _2120_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1140_),
    .A2(net555),
    .Y(_0076_),
    .B1(_0335_));
 sg13g2_o21ai_1 _2121_ (.B1(net625),
    .VDD(VPWR),
    .Y(_0336_),
    .VSS(VGND),
    .A1(net794),
    .A2(net548));
 sg13g2_a21oi_1 _2122_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1139_),
    .A2(net548),
    .Y(_0077_),
    .B1(_0336_));
 sg13g2_o21ai_1 _2123_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0337_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[159] ),
    .A2(net546));
 sg13g2_a21oi_1 _2124_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1138_),
    .A2(net546),
    .Y(_0078_),
    .B1(_0337_));
 sg13g2_o21ai_1 _2125_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0338_),
    .VSS(VGND),
    .A1(net402),
    .A2(net547));
 sg13g2_a21oi_1 _2126_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1137_),
    .A2(net546),
    .Y(_0079_),
    .B1(_0338_));
 sg13g2_o21ai_1 _2127_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0339_),
    .VSS(VGND),
    .A1(net338),
    .A2(net551));
 sg13g2_a21oi_1 _2128_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1136_),
    .A2(net551),
    .Y(_0080_),
    .B1(_0339_));
 sg13g2_o21ai_1 _2129_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0340_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[162] ),
    .A2(net562));
 sg13g2_a21oi_1 _2130_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1135_),
    .A2(net554),
    .Y(_0081_),
    .B1(_0340_));
 sg13g2_o21ai_1 _2131_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0341_),
    .VSS(VGND),
    .A1(net732),
    .A2(net563));
 sg13g2_a21oi_1 _2132_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1134_),
    .A2(net563),
    .Y(_0082_),
    .B1(_0341_));
 sg13g2_o21ai_1 _2133_ (.B1(net633),
    .VDD(VPWR),
    .Y(_0342_),
    .VSS(VGND),
    .A1(net714),
    .A2(net565));
 sg13g2_a21oi_1 _2134_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1133_),
    .A2(net565),
    .Y(_0083_),
    .B1(_0342_));
 sg13g2_o21ai_1 _2135_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0343_),
    .VSS(VGND),
    .A1(net359),
    .A2(net590));
 sg13g2_a21oi_1 _2136_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1132_),
    .A2(net565),
    .Y(_0084_),
    .B1(_0343_));
 sg13g2_o21ai_1 _2137_ (.B1(net655),
    .VDD(VPWR),
    .Y(_0344_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[166] ),
    .A2(net607));
 sg13g2_a21oi_1 _2138_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1131_),
    .A2(net590),
    .Y(_0085_),
    .B1(_0344_));
 sg13g2_o21ai_1 _2139_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0345_),
    .VSS(VGND),
    .A1(net350),
    .A2(net608));
 sg13g2_a21oi_1 _2140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1130_),
    .A2(net608),
    .Y(_0086_),
    .B1(_0345_));
 sg13g2_o21ai_1 _2141_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0346_),
    .VSS(VGND),
    .A1(net336),
    .A2(net616));
 sg13g2_a21oi_1 _2142_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1129_),
    .A2(net608),
    .Y(_0087_),
    .B1(_0346_));
 sg13g2_o21ai_1 _2143_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0347_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[169] ),
    .A2(net615));
 sg13g2_a21oi_1 _2144_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1128_),
    .A2(net615),
    .Y(_0088_),
    .B1(_0347_));
 sg13g2_o21ai_1 _2145_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0348_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[170] ),
    .A2(net619));
 sg13g2_a21oi_1 _2146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1127_),
    .A2(net619),
    .Y(_0089_),
    .B1(_0348_));
 sg13g2_o21ai_1 _2147_ (.B1(net651),
    .VDD(VPWR),
    .Y(_0349_),
    .VSS(VGND),
    .A1(net744),
    .A2(net603));
 sg13g2_a21oi_1 _2148_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1126_),
    .A2(net603),
    .Y(_0090_),
    .B1(_0349_));
 sg13g2_o21ai_1 _2149_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0350_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[172] ),
    .A2(net601));
 sg13g2_a21oi_1 _2150_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1125_),
    .A2(net601),
    .Y(_0091_),
    .B1(_0350_));
 sg13g2_o21ai_1 _2151_ (.B1(net652),
    .VDD(VPWR),
    .Y(_0351_),
    .VSS(VGND),
    .A1(net810),
    .A2(net600));
 sg13g2_a21oi_1 _2152_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1124_),
    .A2(net600),
    .Y(_0092_),
    .B1(_0351_));
 sg13g2_o21ai_1 _2153_ (.B1(net650),
    .VDD(VPWR),
    .Y(_0352_),
    .VSS(VGND),
    .A1(net738),
    .A2(net597));
 sg13g2_a21oi_1 _2154_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1123_),
    .A2(net596),
    .Y(_0093_),
    .B1(_0352_));
 sg13g2_o21ai_1 _2155_ (.B1(net649),
    .VDD(VPWR),
    .Y(_0353_),
    .VSS(VGND),
    .A1(net699),
    .A2(net597));
 sg13g2_a21oi_1 _2156_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1122_),
    .A2(net595),
    .Y(_0094_),
    .B1(_0353_));
 sg13g2_o21ai_1 _2157_ (.B1(net649),
    .VDD(VPWR),
    .Y(_0354_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[176] ),
    .A2(net594));
 sg13g2_a21oi_1 _2158_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1121_),
    .A2(net597),
    .Y(_0095_),
    .B1(_0354_));
 sg13g2_o21ai_1 _2159_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0355_),
    .VSS(VGND),
    .A1(net697),
    .A2(net592));
 sg13g2_a21oi_1 _2160_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1120_),
    .A2(net592),
    .Y(_0096_),
    .B1(_0355_));
 sg13g2_o21ai_1 _2161_ (.B1(net643),
    .VDD(VPWR),
    .Y(_0356_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[178] ),
    .A2(net585));
 sg13g2_a21oi_1 _2162_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1119_),
    .A2(net585),
    .Y(_0097_),
    .B1(_0356_));
 sg13g2_o21ai_1 _2163_ (.B1(net642),
    .VDD(VPWR),
    .Y(_0357_),
    .VSS(VGND),
    .A1(net706),
    .A2(net581));
 sg13g2_a21oi_1 _2164_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1118_),
    .A2(net584),
    .Y(_0098_),
    .B1(_0357_));
 sg13g2_o21ai_1 _2165_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0358_),
    .VSS(VGND),
    .A1(net398),
    .A2(net559));
 sg13g2_a21oi_1 _2166_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1117_),
    .A2(net559),
    .Y(_0099_),
    .B1(_0358_));
 sg13g2_o21ai_1 _2167_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0359_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[181] ),
    .A2(net555));
 sg13g2_a21oi_1 _2168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1116_),
    .A2(net555),
    .Y(_0100_),
    .B1(_0359_));
 sg13g2_o21ai_1 _2169_ (.B1(net625),
    .VDD(VPWR),
    .Y(_0360_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[182] ),
    .A2(net548));
 sg13g2_a21oi_1 _2170_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1115_),
    .A2(net548),
    .Y(_0101_),
    .B1(_0360_));
 sg13g2_o21ai_1 _2171_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0361_),
    .VSS(VGND),
    .A1(net378),
    .A2(net547));
 sg13g2_a21oi_1 _2172_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1114_),
    .A2(net546),
    .Y(_0102_),
    .B1(_0361_));
 sg13g2_o21ai_1 _2173_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0362_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[184] ),
    .A2(net546));
 sg13g2_a21oi_1 _2174_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1113_),
    .A2(net546),
    .Y(_0103_),
    .B1(_0362_));
 sg13g2_o21ai_1 _2175_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0363_),
    .VSS(VGND),
    .A1(net430),
    .A2(net551));
 sg13g2_a21oi_1 _2176_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1112_),
    .A2(net551),
    .Y(_0104_),
    .B1(_0363_));
 sg13g2_o21ai_1 _2177_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0364_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[186] ),
    .A2(net562));
 sg13g2_a21oi_1 _2178_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1111_),
    .A2(net562),
    .Y(_0105_),
    .B1(_0364_));
 sg13g2_o21ai_1 _2179_ (.B1(net634),
    .VDD(VPWR),
    .Y(_0365_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[187] ),
    .A2(net564));
 sg13g2_a21oi_1 _2180_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1110_),
    .A2(net564),
    .Y(_0106_),
    .B1(_0365_));
 sg13g2_o21ai_1 _2181_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0366_),
    .VSS(VGND),
    .A1(net438),
    .A2(net572));
 sg13g2_a21oi_1 _2182_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1109_),
    .A2(net565),
    .Y(_0107_),
    .B1(_0366_));
 sg13g2_o21ai_1 _2183_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0367_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[189] ),
    .A2(net573));
 sg13g2_a21oi_1 _2184_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1108_),
    .A2(net573),
    .Y(_0108_),
    .B1(_0367_));
 sg13g2_o21ai_1 _2185_ (.B1(net655),
    .VDD(VPWR),
    .Y(_0368_),
    .VSS(VGND),
    .A1(net380),
    .A2(net606));
 sg13g2_a21oi_1 _2186_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1107_),
    .A2(net606),
    .Y(_0109_),
    .B1(_0368_));
 sg13g2_o21ai_1 _2187_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0369_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[191] ),
    .A2(net610));
 sg13g2_a21oi_1 _2188_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1106_),
    .A2(net609),
    .Y(_0110_),
    .B1(_0369_));
 sg13g2_o21ai_1 _2189_ (.B1(net662),
    .VDD(VPWR),
    .Y(_0370_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[192] ),
    .A2(net617));
 sg13g2_a21oi_1 _2190_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1105_),
    .A2(net617),
    .Y(_0111_),
    .B1(_0370_));
 sg13g2_o21ai_1 _2191_ (.B1(net662),
    .VDD(VPWR),
    .Y(_0371_),
    .VSS(VGND),
    .A1(net682),
    .A2(net621));
 sg13g2_a21oi_1 _2192_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1104_),
    .A2(net618),
    .Y(_0112_),
    .B1(_0371_));
 sg13g2_o21ai_1 _2193_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0372_),
    .VSS(VGND),
    .A1(net400),
    .A2(net619));
 sg13g2_a21oi_1 _2194_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1103_),
    .A2(net619),
    .Y(_0113_),
    .B1(_0372_));
 sg13g2_o21ai_1 _2195_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0373_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[195] ),
    .A2(net620));
 sg13g2_a21oi_1 _2196_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1102_),
    .A2(net620),
    .Y(_0114_),
    .B1(_0373_));
 sg13g2_o21ai_1 _2197_ (.B1(net651),
    .VDD(VPWR),
    .Y(_0374_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[196] ),
    .A2(net602));
 sg13g2_a21oi_1 _2198_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1101_),
    .A2(net603),
    .Y(_0115_),
    .B1(_0374_));
 sg13g2_o21ai_1 _2199_ (.B1(net652),
    .VDD(VPWR),
    .Y(_0375_),
    .VSS(VGND),
    .A1(net711),
    .A2(net599));
 sg13g2_a21oi_1 _2200_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1100_),
    .A2(net599),
    .Y(_0116_),
    .B1(_0375_));
 sg13g2_o21ai_1 _2201_ (.B1(net652),
    .VDD(VPWR),
    .Y(_0376_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[198] ),
    .A2(net599));
 sg13g2_a21oi_1 _2202_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1099_),
    .A2(net599),
    .Y(_0117_),
    .B1(_0376_));
 sg13g2_o21ai_1 _2203_ (.B1(net649),
    .VDD(VPWR),
    .Y(_0377_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[199] ),
    .A2(net596));
 sg13g2_a21oi_1 _2204_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1098_),
    .A2(net596),
    .Y(_0118_),
    .B1(_0377_));
 sg13g2_o21ai_1 _2205_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0378_),
    .VSS(VGND),
    .A1(\controller.extended_jump_target[0] ),
    .A2(net593));
 sg13g2_a21oi_1 _2206_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1097_),
    .A2(net593),
    .Y(_0119_),
    .B1(_0378_));
 sg13g2_o21ai_1 _2207_ (.B1(net644),
    .VDD(VPWR),
    .Y(_0379_),
    .VSS(VGND),
    .A1(\controller.extended_jump_target[1] ),
    .A2(net587));
 sg13g2_a21oi_1 _2208_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1096_),
    .A2(net587),
    .Y(_0120_),
    .B1(_0379_));
 sg13g2_o21ai_1 _2209_ (.B1(net645),
    .VDD(VPWR),
    .Y(_0380_),
    .VSS(VGND),
    .A1(net842),
    .A2(net583));
 sg13g2_a21oi_1 _2210_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1095_),
    .A2(net583),
    .Y(_0121_),
    .B1(_0380_));
 sg13g2_o21ai_1 _2211_ (.B1(net645),
    .VDD(VPWR),
    .Y(_0381_),
    .VSS(VGND),
    .A1(net729),
    .A2(net582));
 sg13g2_a21oi_1 _2212_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1094_),
    .A2(net582),
    .Y(_0122_),
    .B1(_0381_));
 sg13g2_o21ai_1 _2213_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0382_),
    .VSS(VGND),
    .A1(net334),
    .A2(net561));
 sg13g2_a21oi_1 _2214_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1093_),
    .A2(net561),
    .Y(_0123_),
    .B1(_0382_));
 sg13g2_o21ai_1 _2215_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0383_),
    .VSS(VGND),
    .A1(\controller.inst_mem.extended_word[5] ),
    .A2(net556));
 sg13g2_a21oi_1 _2216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1092_),
    .A2(net561),
    .Y(_0124_),
    .B1(_0383_));
 sg13g2_o21ai_1 _2217_ (.B1(net628),
    .VDD(VPWR),
    .Y(_0384_),
    .VSS(VGND),
    .A1(net701),
    .A2(net557));
 sg13g2_a21oi_1 _2218_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1091_),
    .A2(net557),
    .Y(_0125_),
    .B1(_0384_));
 sg13g2_o21ai_1 _2219_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0385_),
    .VSS(VGND),
    .A1(\controller.inst_mem.extended_word[7] ),
    .A2(net549));
 sg13g2_a21oi_1 _2220_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1090_),
    .A2(net549),
    .Y(_0126_),
    .B1(_0385_));
 sg13g2_o21ai_1 _2221_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0386_),
    .VSS(VGND),
    .A1(net761),
    .A2(net551));
 sg13g2_a21oi_1 _2222_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1089_),
    .A2(net551),
    .Y(_0127_),
    .B1(_0386_));
 sg13g2_o21ai_1 _2223_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0387_),
    .VSS(VGND),
    .A1(\controller.extended_cond.opcode[0] ),
    .A2(net554));
 sg13g2_a21oi_1 _2224_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1088_),
    .A2(net554),
    .Y(_0128_),
    .B1(_0387_));
 sg13g2_o21ai_1 _2225_ (.B1(net639),
    .VDD(VPWR),
    .Y(_0388_),
    .VSS(VGND),
    .A1(\controller.extended_cond.opcode[1] ),
    .A2(net575));
 sg13g2_a21oi_1 _2226_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1087_),
    .A2(net575),
    .Y(_0129_),
    .B1(_0388_));
 sg13g2_o21ai_1 _2227_ (.B1(net639),
    .VDD(VPWR),
    .Y(_0389_),
    .VSS(VGND),
    .A1(net885),
    .A2(net575));
 sg13g2_a21oi_1 _2228_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1086_),
    .A2(net575),
    .Y(_0130_),
    .B1(_0389_));
 sg13g2_o21ai_1 _2229_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0390_),
    .VSS(VGND),
    .A1(net858),
    .A2(net575));
 sg13g2_a21oi_1 _2230_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1085_),
    .A2(net575),
    .Y(_0131_),
    .B1(_0390_));
 sg13g2_o21ai_1 _2231_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0391_),
    .VSS(VGND),
    .A1(net728),
    .A2(net572));
 sg13g2_a21oi_1 _2232_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1084_),
    .A2(net572),
    .Y(_0132_),
    .B1(_0391_));
 sg13g2_o21ai_1 _2233_ (.B1(net655),
    .VDD(VPWR),
    .Y(_0392_),
    .VSS(VGND),
    .A1(net685),
    .A2(net607));
 sg13g2_a21oi_1 _2234_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1083_),
    .A2(net607),
    .Y(_0133_),
    .B1(_0392_));
 sg13g2_o21ai_1 _2235_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(\controller.extended_then_action[3] ),
    .A2(net608));
 sg13g2_a21oi_1 _2236_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1082_),
    .A2(net608),
    .Y(_0134_),
    .B1(_0393_));
 sg13g2_o21ai_1 _2237_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0394_),
    .VSS(VGND),
    .A1(net881),
    .A2(net611));
 sg13g2_a21oi_1 _2238_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1081_),
    .A2(net611),
    .Y(_0135_),
    .B1(_0394_));
 sg13g2_o21ai_1 _2239_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0395_),
    .VSS(VGND),
    .A1(net878),
    .A2(net616));
 sg13g2_a21oi_1 _2240_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1080_),
    .A2(net616),
    .Y(_0136_),
    .B1(_0395_));
 sg13g2_o21ai_1 _2241_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0396_),
    .VSS(VGND),
    .A1(net364),
    .A2(net615));
 sg13g2_a21oi_1 _2242_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1079_),
    .A2(net615),
    .Y(_0137_),
    .B1(_0396_));
 sg13g2_o21ai_1 _2243_ (.B1(net651),
    .VDD(VPWR),
    .Y(_0397_),
    .VSS(VGND),
    .A1(\controller.inst_mem.extended_word[19] ),
    .A2(net602));
 sg13g2_a21oi_1 _2244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1078_),
    .A2(net602),
    .Y(_0138_),
    .B1(_0397_));
 sg13g2_o21ai_1 _2245_ (.B1(net651),
    .VDD(VPWR),
    .Y(_0398_),
    .VSS(VGND),
    .A1(\controller.inst_mem.extended_word[20] ),
    .A2(net602));
 sg13g2_a21oi_1 _2246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1077_),
    .A2(net602),
    .Y(_0139_),
    .B1(_0398_));
 sg13g2_o21ai_1 _2247_ (.B1(net652),
    .VDD(VPWR),
    .Y(_0399_),
    .VSS(VGND),
    .A1(\controller.inst_mem.extended_word[21] ),
    .A2(net599));
 sg13g2_a21oi_1 _2248_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1076_),
    .A2(net599),
    .Y(_0140_),
    .B1(_0399_));
 sg13g2_o21ai_1 _2249_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0400_),
    .VSS(VGND),
    .A1(net353),
    .A2(net598));
 sg13g2_a21oi_1 _2250_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1075_),
    .A2(net598),
    .Y(_0141_),
    .B1(_0400_));
 sg13g2_o21ai_1 _2251_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0401_),
    .VSS(VGND),
    .A1(\controller.inst_mem.extended_word[23] ),
    .A2(net593));
 sg13g2_a21oi_1 _2252_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1074_),
    .A2(net598),
    .Y(_0142_),
    .B1(_0401_));
 sg13g2_o21ai_1 _2253_ (.B1(net647),
    .VDD(VPWR),
    .Y(_0402_),
    .VSS(VGND),
    .A1(net376),
    .A2(net589));
 sg13g2_a21oi_1 _2254_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1073_),
    .A2(net589),
    .Y(_0143_),
    .B1(_0402_));
 sg13g2_o21ai_1 _2255_ (.B1(net647),
    .VDD(VPWR),
    .Y(_0403_),
    .VSS(VGND),
    .A1(\controller.extended_state[1] ),
    .A2(net589));
 sg13g2_a21oi_1 _2256_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1072_),
    .A2(net589),
    .Y(_0144_),
    .B1(_0403_));
 sg13g2_o21ai_1 _2257_ (.B1(net647),
    .VDD(VPWR),
    .Y(_0404_),
    .VSS(VGND),
    .A1(\controller.extended_state[2] ),
    .A2(net588));
 sg13g2_a21oi_1 _2258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1071_),
    .A2(net588),
    .Y(_0145_),
    .B1(_0404_));
 sg13g2_nor2_1 _2259_ (.A(net930),
    .B(\controller.counter2.counter_0[0] ),
    .Y(_0405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2260_ (.A(net919),
    .B(\controller.counter2.counter_0[1] ),
    .C(\controller.counter2.counter_0[0] ),
    .Y(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _2261_ (.A(\controller.counter2.counter_0[3] ),
    .B(\controller.counter2.counter_0[2] ),
    .C(\controller.counter2.counter_0[1] ),
    .D(\controller.counter2.counter_0[0] ),
    .X(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2262_ (.A(net944),
    .B(_0407_),
    .Y(_0408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2263_ (.A(net938),
    .B(\controller.counter2.counter_0[4] ),
    .C(_0407_),
    .Y(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2264_ (.A(net894),
    .B(\controller.counter2.counter_0[5] ),
    .C(\controller.counter2.counter_0[4] ),
    .Y(_0410_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0407_));
 sg13g2_nand2_1 _2265_ (.Y(_0411_),
    .A(_1063_),
    .B(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2266_ (.A(\controller.counter2.counter_0[9] ),
    .B(\controller.counter2.counter_0[8] ),
    .Y(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2267_ (.B(_0410_),
    .C(_0412_),
    .A(_1063_),
    .Y(_0413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2268_ (.B(_1063_),
    .C(_0410_),
    .A(_1062_),
    .Y(_0414_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0412_));
 sg13g2_or2_1 _2269_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0415_),
    .B(_0414_),
    .A(net897));
 sg13g2_or2_1 _2270_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0416_),
    .B(\controller.counter2.counter_0[12] ),
    .A(\controller.counter2.counter_0[13] ));
 sg13g2_nor2_1 _2271_ (.A(_0415_),
    .B(_0416_),
    .Y(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2272_ (.A(net893),
    .B(net897),
    .C(_0414_),
    .D(_0416_),
    .Y(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2273_ (.Y(_0419_),
    .B(_0418_),
    .A_N(\controller.counter2.counter_0[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2274_ (.A(\controller.extended_cond.opcode[2] ),
    .B(\controller.extended_cond.opcode[1] ),
    .Y(_0420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2275_ (.A(\controller.extended_cond.opcode[2] ),
    .B(\controller.extended_cond.opcode[1] ),
    .C(\controller.extended_cond.opcode[0] ),
    .Y(_0421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2276_ (.A(_0419_),
    .B(_0421_),
    .X(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2277_ (.B(\controller.extended_state[2] ),
    .A(net532),
    .X(_0423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2278_ (.B(\controller.extended_state[1] ),
    .A(net534),
    .X(_0424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2279_ (.B(\controller.extended_state[0] ),
    .A(net535),
    .X(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2280_ (.A(net524),
    .B(_0423_),
    .C(_0424_),
    .D(_0425_),
    .Y(_0426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2281_ (.Y(_0427_),
    .A(\controller.extended_cond.opcode[2] ),
    .B(\controller.extended_cond.opcode[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2282_ (.A(net2),
    .B(_0427_),
    .Y(_0428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2283_ (.B1(_1086_),
    .VDD(VPWR),
    .Y(_0429_),
    .VSS(VGND),
    .A1(\controller.extended_cond.opcode[0] ),
    .A2(net1));
 sg13g2_nand2_1 _2284_ (.Y(_0430_),
    .A(_1085_),
    .B(\controller.extended_cond.opcode[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2285_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0429_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(_0428_));
 sg13g2_nor2_1 _2286_ (.A(net4),
    .B(_0427_),
    .Y(_0432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2287_ (.B1(\controller.extended_cond.opcode[1] ),
    .VDD(VPWR),
    .Y(_0433_),
    .VSS(VGND),
    .A1(\controller.extended_cond.opcode[0] ),
    .A2(net3));
 sg13g2_nor2_1 _2288_ (.A(_0432_),
    .B(_0433_),
    .Y(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2289_ (.A(_0431_),
    .B(_0434_),
    .Y(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2290_ (.A(_1087_),
    .B(_0430_),
    .Y(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2291_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1300_),
    .C1(_0435_),
    .B1(_0436_),
    .A1(_1280_),
    .Y(_0437_),
    .A2(_0420_));
 sg13g2_o21ai_1 _2292_ (.B1(_0426_),
    .VDD(VPWR),
    .Y(_0438_),
    .VSS(VGND),
    .A1(_0421_),
    .A2(_0437_));
 sg13g2_or2_1 _2293_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0439_),
    .B(net489),
    .A(_0422_));
 sg13g2_nor2_1 _2294_ (.A(net844),
    .B(net488),
    .Y(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2295_ (.A(_1110_),
    .B(_1223_),
    .Y(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2296_ (.B(net533),
    .C(net536),
    .A(net532),
    .Y(_0442_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\controller.extended_cond.opcode[1] ));
 sg13g2_nor3_1 _2297_ (.A(net531),
    .B(_1206_),
    .C(_1221_),
    .Y(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2298_ (.A(\controller.inst_mem.mem_data[138] ),
    .B(net519),
    .X(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2299_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[114] ),
    .C1(_0443_),
    .B1(net498),
    .A1(\controller.inst_mem.mem_data[66] ),
    .Y(_0445_),
    .A2(net509));
 sg13g2_o21ai_1 _2300_ (.B1(_0442_),
    .VDD(VPWR),
    .Y(_0446_),
    .VSS(VGND),
    .A1(_1134_),
    .A2(_1218_));
 sg13g2_nor4_1 _2301_ (.A(net515),
    .B(_0441_),
    .C(_0444_),
    .D(_0446_),
    .Y(_0447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2302_ (.Y(_0448_),
    .B1(_0445_),
    .B2(_0447_),
    .A2(net515),
    .A1(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2303_ (.A(\controller.extended_cond.opcode[2] ),
    .B(net523),
    .X(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2304_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[67] ),
    .C1(_0449_),
    .B1(net506),
    .A1(\controller.inst_mem.mem_data[163] ),
    .Y(_0450_),
    .A2(net510));
 sg13g2_nor3_1 _2305_ (.A(net531),
    .B(_1205_),
    .C(_1221_),
    .Y(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2306_ (.A2(net519),
    .A1(\controller.inst_mem.mem_data[139] ),
    .B1(net515),
    .X(_0452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2307_ (.A(net531),
    .B(_1181_),
    .C(_1225_),
    .Y(_0453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2308_ (.A(_1109_),
    .B(_1223_),
    .Y(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2309_ (.A(_0451_),
    .B(_0452_),
    .C(_0453_),
    .D(_0454_),
    .Y(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2310_ (.A(\controller.inst_mem.mem_data[43] ),
    .B(net493),
    .Y(_0456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _2311_ (.A2(_0455_),
    .A1(_0450_),
    .B1(_0456_),
    .X(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2312_ (.A(_0448_),
    .B_N(_0457_),
    .Y(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2313_ (.Y(_0459_),
    .A(\controller.inst_mem.mem_data[89] ),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2314_ (.Y(_0460_),
    .B1(net523),
    .B2(\controller.extended_cond.opcode[0] ),
    .A2(net506),
    .A1(\controller.inst_mem.mem_data[65] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2315_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[137] ),
    .C1(net514),
    .B1(net519),
    .A1(\controller.inst_mem.mem_data[113] ),
    .Y(_0461_),
    .A2(net498));
 sg13g2_a22oi_1 _2316_ (.Y(_0462_),
    .B1(net502),
    .B2(\controller.inst_mem.mem_data[185] ),
    .A2(net510),
    .A1(\controller.inst_mem.mem_data[161] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2317_ (.B(_0460_),
    .C(_0461_),
    .A(_0459_),
    .Y(_0463_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0462_));
 sg13g2_nand2_1 _2318_ (.Y(_0464_),
    .A(_1019_),
    .B(net515),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2319_ (.A(_0463_),
    .B(_0464_),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2320_ (.Y(_0466_),
    .A(_0463_),
    .B(_0464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2321_ (.Y(_0467_),
    .B(net1),
    .A_N(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2322_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3),
    .A2(_0448_),
    .Y(_0468_),
    .B1(_0457_));
 sg13g2_a221oi_1 _2323_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0468_),
    .C1(_0465_),
    .B1(_0467_),
    .A1(_0419_),
    .Y(_0469_),
    .A2(_0458_));
 sg13g2_mux2_1 _2324_ (.A0(_1280_),
    .A1(_1300_),
    .S(_0448_),
    .X(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2325_ (.Y(_0471_),
    .B(net2),
    .A_N(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2326_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net4),
    .A2(_0448_),
    .Y(_0472_),
    .B1(_0457_));
 sg13g2_a221oi_1 _2327_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0472_),
    .C1(_0466_),
    .B1(_0471_),
    .A1(_0457_),
    .Y(_0473_),
    .A2(_0470_));
 sg13g2_nor2_1 _2328_ (.A(_0469_),
    .B(_0473_),
    .Y(_0474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2329_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0475_),
    .B(_0473_),
    .A(_0469_));
 sg13g2_a21oi_1 _2330_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net535),
    .A2(net488),
    .Y(_0476_),
    .B1(_0440_));
 sg13g2_nand2_1 _2331_ (.Y(_0477_),
    .A(net486),
    .B(_0476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2332_ (.Y(_0478_),
    .B1(net494),
    .B2(\controller.inst_mem.mem_data[84] ),
    .A2(net506),
    .A1(\controller.inst_mem.mem_data[60] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2333_ (.A(net532),
    .B(net522),
    .X(_0479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2334_ (.Y(_0480_),
    .B1(net502),
    .B2(\controller.inst_mem.mem_data[180] ),
    .A2(net510),
    .A1(\controller.inst_mem.mem_data[156] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2335_ (.Y(_0481_),
    .B1(_0479_),
    .B2(\controller.inst_mem.mem_data[132] ),
    .A2(net523),
    .A1(\controller.inst_mem.extended_word[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2336_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[108] ),
    .A2(net498),
    .Y(_0482_),
    .B1(net516));
 sg13g2_nand4_1 _2337_ (.B(_0480_),
    .C(_0481_),
    .A(_0478_),
    .Y(_0483_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0482_));
 sg13g2_nand2_1 _2338_ (.Y(_0484_),
    .A(_1280_),
    .B(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2339_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0484_),
    .Y(_0485_),
    .A2(net515),
    .A1(_1024_));
 sg13g2_a21o_2 _2340_ (.A2(net515),
    .A1(_1024_),
    .B1(_0484_),
    .X(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2341_ (.Y(_0487_),
    .B1(net523),
    .B2(\controller.inst_mem.extended_word[3] ),
    .A2(net506),
    .A1(\controller.inst_mem.mem_data[59] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2342_ (.Y(_0488_),
    .A(\controller.inst_mem.mem_data[179] ),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2343_ (.Y(_0489_),
    .B1(net494),
    .B2(\controller.inst_mem.mem_data[83] ),
    .A2(net510),
    .A1(\controller.inst_mem.mem_data[155] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2344_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[131] ),
    .C1(net517),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[107] ),
    .Y(_0490_),
    .A2(net498));
 sg13g2_nand4_1 _2345_ (.B(_0488_),
    .C(_0489_),
    .A(_0487_),
    .Y(_0491_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0490_));
 sg13g2_nand2_1 _2346_ (.Y(_0492_),
    .A(_1025_),
    .B(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2347_ (.B(net486),
    .C(_0491_),
    .A(net488),
    .Y(_0493_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0492_));
 sg13g2_nand2_2 _2348_ (.Y(_0494_),
    .A(_0486_),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2349_ (.Y(_0495_),
    .B1(net524),
    .B2(\controller.extended_jump_target[0] ),
    .A2(net499),
    .A1(\controller.inst_mem.mem_data[104] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2350_ (.Y(_0496_),
    .B1(net495),
    .B2(\controller.inst_mem.mem_data[80] ),
    .A2(net507),
    .A1(\controller.inst_mem.mem_data[56] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2351_ (.Y(_0497_),
    .B1(_0479_),
    .B2(\controller.inst_mem.mem_data[128] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[152] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2352_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[176] ),
    .A2(net503),
    .Y(_0498_),
    .B1(net517));
 sg13g2_nand4_1 _2353_ (.B(_0496_),
    .C(_0497_),
    .A(_0495_),
    .Y(_0499_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0498_));
 sg13g2_o21ai_1 _2354_ (.B1(_0499_),
    .VDD(VPWR),
    .Y(_0500_),
    .VSS(VGND),
    .A1(net777),
    .A2(net491));
 sg13g2_o21ai_1 _2355_ (.B1(_0477_),
    .VDD(VPWR),
    .Y(_0501_),
    .VSS(VGND),
    .A1(net486),
    .A2(_0500_));
 sg13g2_nor2b_2 _2356_ (.A(net6),
    .B_N(net637),
    .Y(_0502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2357_ (.Y(_0503_),
    .B(net637),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net6));
 sg13g2_o21ai_1 _2358_ (.B1(net545),
    .VDD(VPWR),
    .Y(_0504_),
    .VSS(VGND),
    .A1(_0494_),
    .A2(_0501_));
 sg13g2_a21oi_1 _2359_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1070_),
    .A2(_0494_),
    .Y(_0146_),
    .B1(_0504_));
 sg13g2_xnor2_1 _2360_ (.Y(_0505_),
    .A(net534),
    .B(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[57] ),
    .A2(net507),
    .Y(_0506_),
    .B1(net517));
 sg13g2_a22oi_1 _2362_ (.Y(_0507_),
    .B1(net495),
    .B2(\controller.inst_mem.mem_data[81] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[153] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2363_ (.Y(_0508_),
    .B1(net499),
    .B2(\controller.inst_mem.mem_data[105] ),
    .A2(net503),
    .A1(\controller.inst_mem.mem_data[177] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2364_ (.Y(_0509_),
    .B1(_0479_),
    .B2(\controller.inst_mem.mem_data[129] ),
    .A2(net524),
    .A1(\controller.extended_jump_target[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2365_ (.B(_0507_),
    .C(_0508_),
    .A(_0506_),
    .Y(_0510_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0509_));
 sg13g2_o21ai_1 _2366_ (.B1(_0510_),
    .VDD(VPWR),
    .Y(_0511_),
    .VSS(VGND),
    .A1(net720),
    .A2(net491));
 sg13g2_o21ai_1 _2367_ (.B1(net486),
    .VDD(VPWR),
    .Y(_0512_),
    .VSS(VGND),
    .A1(net854),
    .A2(net488));
 sg13g2_a21o_1 _2368_ (.A2(_0505_),
    .A1(net488),
    .B1(_0512_),
    .X(_0513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2369_ (.A(net486),
    .B(_0511_),
    .Y(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2370_ (.A(_0494_),
    .B(_0514_),
    .Y(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2371_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0515_),
    .C1(_0503_),
    .B1(_0513_),
    .A1(_1069_),
    .Y(_0147_),
    .A2(_0494_));
 sg13g2_a21oi_1 _2372_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net534),
    .A2(net535),
    .Y(_0516_),
    .B1(net531));
 sg13g2_o21ai_1 _2373_ (.B1(net488),
    .VDD(VPWR),
    .Y(_0517_),
    .VSS(VGND),
    .A1(net524),
    .A2(_0516_));
 sg13g2_a22oi_1 _2374_ (.Y(_0518_),
    .B1(net524),
    .B2(\controller.extended_jump_target[2] ),
    .A2(net507),
    .A1(\controller.inst_mem.mem_data[58] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2375_ (.Y(_0519_),
    .B1(net499),
    .B2(\controller.inst_mem.mem_data[106] ),
    .A2(net503),
    .A1(\controller.inst_mem.mem_data[178] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2376_ (.Y(_0520_),
    .B1(_0479_),
    .B2(\controller.inst_mem.mem_data[130] ),
    .A2(net495),
    .A1(\controller.inst_mem.mem_data[82] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2377_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[154] ),
    .A2(net511),
    .Y(_0521_),
    .B1(net517));
 sg13g2_nand4_1 _2378_ (.B(_0519_),
    .C(_0520_),
    .A(_0518_),
    .Y(_0522_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0521_));
 sg13g2_o21ai_1 _2379_ (.B1(_0522_),
    .VDD(VPWR),
    .Y(_0523_),
    .VSS(VGND),
    .A1(net800),
    .A2(net491));
 sg13g2_o21ai_1 _2380_ (.B1(net486),
    .VDD(VPWR),
    .Y(_0524_),
    .VSS(VGND),
    .A1(\controller.extended_jump_target[2] ),
    .A2(net488));
 sg13g2_nand2b_1 _2381_ (.Y(_0525_),
    .B(_0517_),
    .A_N(_0524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2382_ (.B1(_0525_),
    .VDD(VPWR),
    .Y(_0526_),
    .VSS(VGND),
    .A1(net486),
    .A2(_0523_));
 sg13g2_o21ai_1 _2383_ (.B1(net545),
    .VDD(VPWR),
    .Y(_0527_),
    .VSS(VGND),
    .A1(_0494_),
    .A2(_0526_));
 sg13g2_a21oi_1 _2384_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1068_),
    .A2(_0494_),
    .Y(_0148_),
    .B1(_0527_));
 sg13g2_or3_1 _2385_ (.A(_1080_),
    .B(net490),
    .C(net489),
    .X(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2386_ (.Y(_0529_),
    .A(\controller.inst_mem.extended_word[22] ),
    .B(net524),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2387_ (.Y(_0530_),
    .B1(net499),
    .B2(\controller.inst_mem.mem_data[126] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[174] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2388_ (.Y(_0531_),
    .B1(net503),
    .B2(\controller.inst_mem.mem_data[198] ),
    .A2(net507),
    .A1(\controller.inst_mem.mem_data[78] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2389_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[150] ),
    .C1(net517),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[102] ),
    .Y(_0532_),
    .A2(net495));
 sg13g2_nand4_1 _2390_ (.B(_0530_),
    .C(_0531_),
    .A(_0529_),
    .Y(_0533_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0532_));
 sg13g2_o21ai_1 _2391_ (.B1(_0533_),
    .VDD(VPWR),
    .Y(_0534_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[54] ),
    .A2(net491));
 sg13g2_inv_1 _2392_ (.VDD(VPWR),
    .Y(_0535_),
    .A(_0534_),
    .VSS(VGND));
 sg13g2_o21ai_1 _2393_ (.B1(_0535_),
    .VDD(VPWR),
    .Y(_0536_),
    .VSS(VGND),
    .A1(net490),
    .A2(net489));
 sg13g2_nand3_1 _2394_ (.B(_0528_),
    .C(_0536_),
    .A(net486),
    .Y(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2395_ (.Y(_0538_),
    .A(\controller.inst_mem.mem_data[120] ),
    .B(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2396_ (.Y(_0539_),
    .B1(net495),
    .B2(\controller.inst_mem.mem_data[96] ),
    .A2(net503),
    .A1(\controller.inst_mem.mem_data[192] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2397_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[144] ),
    .C1(net518),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[72] ),
    .Y(_0540_),
    .A2(net507));
 sg13g2_a22oi_1 _2398_ (.Y(_0541_),
    .B1(net525),
    .B2(\controller.extended_then_action[4] ),
    .A2(net512),
    .A1(\controller.inst_mem.mem_data[168] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2399_ (.B(_0539_),
    .C(_0540_),
    .A(_0538_),
    .Y(_0542_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0541_));
 sg13g2_o21ai_1 _2400_ (.B1(_0542_),
    .VDD(VPWR),
    .Y(_0543_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[48] ),
    .A2(net492));
 sg13g2_a21oi_1 _2401_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0543_),
    .Y(_0544_),
    .B1(_0485_));
 sg13g2_and2_1 _2402_ (.A(_0537_),
    .B(_0544_),
    .X(_0545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2403_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0546_),
    .B(_0439_),
    .A(_1079_));
 sg13g2_a221oi_1 _2404_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[151] ),
    .C1(net518),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[127] ),
    .Y(_0547_),
    .A2(net499));
 sg13g2_a22oi_1 _2405_ (.Y(_0548_),
    .B1(net495),
    .B2(\controller.inst_mem.mem_data[103] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[175] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2406_ (.Y(_0549_),
    .B1(net503),
    .B2(\controller.inst_mem.mem_data[199] ),
    .A2(net507),
    .A1(\controller.inst_mem.mem_data[79] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2407_ (.B(_0548_),
    .C(_0549_),
    .A(_0547_),
    .Y(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2408_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.extended_word[23] ),
    .A2(net524),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_a21oi_2 _2409_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0551_),
    .Y(_0552_),
    .A2(net517),
    .A1(_1005_));
 sg13g2_a21oi_1 _2410_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0439_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(_0475_));
 sg13g2_nand2_1 _2411_ (.Y(_0554_),
    .A(\controller.inst_mem.mem_data[121] ),
    .B(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2412_ (.Y(_0555_),
    .B1(net503),
    .B2(\controller.inst_mem.mem_data[193] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[169] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2413_ (.Y(_0556_),
    .B1(net525),
    .B2(\controller.extended_then_action[5] ),
    .A2(net507),
    .A1(\controller.inst_mem.mem_data[73] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2414_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[145] ),
    .C1(net518),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[97] ),
    .Y(_0557_),
    .A2(net495));
 sg13g2_nand4_1 _2415_ (.B(_0555_),
    .C(_0556_),
    .A(_0554_),
    .Y(_0558_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0557_));
 sg13g2_o21ai_1 _2416_ (.B1(_0558_),
    .VDD(VPWR),
    .Y(_0559_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[49] ),
    .A2(net491));
 sg13g2_a21o_1 _2417_ (.A2(_0559_),
    .A1(_0475_),
    .B1(_0485_),
    .X(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2418_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0560_),
    .Y(_0561_),
    .A2(_0553_),
    .A1(_0546_));
 sg13g2_or2_1 _2419_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0562_),
    .B(_0561_),
    .A(net485));
 sg13g2_nor2_1 _2420_ (.A(\controller.alu_buffer.buffer[0] ),
    .B(_0562_),
    .Y(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2421_ (.A(_1081_),
    .B(net490),
    .C(_0438_),
    .X(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2422_ (.Y(_0565_),
    .A(\controller.inst_mem.mem_data[197] ),
    .B(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2423_ (.Y(_0566_),
    .B1(net524),
    .B2(\controller.inst_mem.extended_word[21] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[173] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2424_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[149] ),
    .C1(net517),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[125] ),
    .Y(_0567_),
    .A2(net499));
 sg13g2_a22oi_1 _2425_ (.Y(_0568_),
    .B1(net495),
    .B2(\controller.inst_mem.mem_data[101] ),
    .A2(net507),
    .A1(\controller.inst_mem.mem_data[77] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2426_ (.B(_0566_),
    .C(_0567_),
    .A(_0565_),
    .Y(_0569_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0568_));
 sg13g2_o21ai_1 _2427_ (.B1(_0569_),
    .VDD(VPWR),
    .Y(_0570_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[53] ),
    .A2(net491));
 sg13g2_inv_1 _2428_ (.VDD(VPWR),
    .Y(_0571_),
    .A(_0570_),
    .VSS(VGND));
 sg13g2_o21ai_1 _2429_ (.B1(_0571_),
    .VDD(VPWR),
    .Y(_0572_),
    .VSS(VGND),
    .A1(net490),
    .A2(net489));
 sg13g2_nand3_1 _2430_ (.B(_0564_),
    .C(_0572_),
    .A(net487),
    .Y(_0573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2431_ (.Y(_0574_),
    .A(\controller.inst_mem.mem_data[71] ),
    .B(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2432_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[143] ),
    .C1(net518),
    .B1(net520),
    .A1(\controller.inst_mem.mem_data[167] ),
    .Y(_0575_),
    .A2(net512));
 sg13g2_a22oi_1 _2433_ (.Y(_0576_),
    .B1(net525),
    .B2(\controller.extended_then_action[3] ),
    .A2(net500),
    .A1(\controller.inst_mem.mem_data[119] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2434_ (.Y(_0577_),
    .B1(net496),
    .B2(\controller.inst_mem.mem_data[95] ),
    .A2(net504),
    .A1(\controller.inst_mem.mem_data[191] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2435_ (.B(_0575_),
    .C(_0576_),
    .A(_0574_),
    .Y(_0578_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0577_));
 sg13g2_o21ai_1 _2436_ (.B1(_0578_),
    .VDD(VPWR),
    .Y(_0579_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[47] ),
    .A2(net492));
 sg13g2_a21oi_1 _2437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(_0485_));
 sg13g2_and2_1 _2438_ (.A(_0573_),
    .B(_0580_),
    .X(_0581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2439_ (.Y(_0582_),
    .A(_0573_),
    .B(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2440_ (.Y(_0583_),
    .A(net485),
    .B(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2441_ (.X(_0584_),
    .A(net485),
    .B(_0561_),
    .C(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2442_ (.Y(_0585_),
    .A(\controller.alu_buffer.buffer[7] ),
    .B(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2443_ (.X(_0586_),
    .A(net485),
    .B(_0561_),
    .C(_0581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2444_ (.Y(_0587_),
    .A(\controller.alu_buffer.buffer[8] ),
    .B(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2445_ (.B(net527),
    .A(\controller.alu_buffer.buffer[7] ),
    .X(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2446_ (.B(net528),
    .A(\controller.alu_buffer.buffer[5] ),
    .X(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2447_ (.Y(_0590_),
    .A(_0588_),
    .B(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2448_ (.Y(_0591_),
    .A(net530),
    .B(net971),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2449_ (.B(net529),
    .A(\controller.alu_buffer.buffer[3] ),
    .X(_0592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2450_ (.Y(_0593_),
    .A(_0591_),
    .B(_0592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2451_ (.Y(_0594_),
    .A(_0590_),
    .B(_0593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2452_ (.A(_0561_),
    .B(_0581_),
    .Y(_0595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2453_ (.Y(_0596_),
    .B(_0582_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0561_));
 sg13g2_and2_1 _2454_ (.A(net485),
    .B(_0594_),
    .X(_0597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1065_),
    .A2(_0561_),
    .Y(_0598_),
    .B1(net485));
 sg13g2_a221oi_1 _2456_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0597_),
    .C1(_0598_),
    .B1(net463),
    .A1(net468),
    .Y(_0599_),
    .A2(_0587_));
 sg13g2_a21o_1 _2457_ (.A2(_0599_),
    .A1(_0585_),
    .B1(_0563_),
    .X(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2458_ (.Y(_0601_),
    .B(net463),
    .A_N(_0545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2459_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0602_),
    .VSS(VGND),
    .A1(net967),
    .A2(_0601_));
 sg13g2_a21oi_1 _2460_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0600_),
    .A2(_0601_),
    .Y(_0149_),
    .B1(_0602_));
 sg13g2_a221oi_1 _2461_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0553_),
    .C1(_0560_),
    .B1(_0546_),
    .A1(_0537_),
    .Y(_0603_),
    .A2(_0544_));
 sg13g2_a22oi_1 _2462_ (.Y(_0604_),
    .B1(net460),
    .B2(_1061_),
    .A2(_0583_),
    .A1(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2463_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net530),
    .C1(_0604_),
    .B1(net484),
    .A1(_1067_),
    .Y(_0605_),
    .A2(net468));
 sg13g2_o21ai_1 _2464_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0606_),
    .VSS(VGND),
    .A1(net971),
    .A2(_0596_));
 sg13g2_nor2_1 _2465_ (.A(_0605_),
    .B(_0606_),
    .Y(_0150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2466_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0561_),
    .Y(_0607_),
    .A2(_0581_),
    .A1(net485));
 sg13g2_a22oi_1 _2467_ (.Y(_0608_),
    .B1(net457),
    .B2(net8),
    .A2(_0591_),
    .A1(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2468_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net529),
    .C1(net463),
    .B1(net483),
    .A1(net971),
    .Y(_0609_),
    .A2(net473));
 sg13g2_o21ai_1 _2469_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0610_),
    .VSS(VGND),
    .A1(net530),
    .A2(net460));
 sg13g2_a21oi_1 _2470_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0608_),
    .A2(_0609_),
    .Y(_0151_),
    .B1(_0610_));
 sg13g2_a221oi_1 _2471_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net977),
    .C1(net463),
    .B1(net483),
    .A1(net530),
    .Y(_0611_),
    .A2(net472));
 sg13g2_or3_1 _2472_ (.A(net529),
    .B(net530),
    .C(net984),
    .X(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2473_ (.B1(net529),
    .VDD(VPWR),
    .Y(_0613_),
    .VSS(VGND),
    .A1(net530),
    .A2(net984));
 sg13g2_nand2_1 _2474_ (.Y(_0614_),
    .A(_0612_),
    .B(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2475_ (.Y(_0615_),
    .B1(_0614_),
    .B2(net468),
    .A2(net457),
    .A1(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2476_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0616_),
    .VSS(VGND),
    .A1(net529),
    .A2(net460));
 sg13g2_a21oi_1 _2477_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0611_),
    .A2(_0615_),
    .Y(_0152_),
    .B1(_0616_));
 sg13g2_a21o_1 _2478_ (.A2(_0612_),
    .A1(net977),
    .B1(_1283_),
    .X(_0617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2479_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net468),
    .C1(net463),
    .B1(_0617_),
    .A1(net528),
    .Y(_0618_),
    .A2(net483));
 sg13g2_a22oi_1 _2480_ (.Y(_0619_),
    .B1(net457),
    .B2(net10),
    .A2(net472),
    .A1(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2481_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0620_),
    .VSS(VGND),
    .A1(net977),
    .A2(net460));
 sg13g2_a21oi_1 _2482_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0618_),
    .A2(_0619_),
    .Y(_0153_),
    .B1(_0620_));
 sg13g2_a221oi_1 _2483_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net980),
    .C1(net463),
    .B1(net483),
    .A1(net977),
    .Y(_0621_),
    .A2(net472));
 sg13g2_nor2b_1 _2484_ (.A(net528),
    .B_N(_1283_),
    .Y(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2485_ (.B(_1283_),
    .A(net528),
    .X(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2486_ (.Y(_0624_),
    .B1(_0623_),
    .B2(net468),
    .A2(net457),
    .A1(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2487_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0625_),
    .VSS(VGND),
    .A1(net528),
    .A2(net460));
 sg13g2_a21oi_1 _2488_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0621_),
    .A2(_0624_),
    .Y(_0154_),
    .B1(_0625_));
 sg13g2_o21ai_1 _2489_ (.B1(_1285_),
    .VDD(VPWR),
    .Y(_0626_),
    .VSS(VGND),
    .A1(_1066_),
    .A2(_0622_));
 sg13g2_a221oi_1 _2490_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net469),
    .C1(net464),
    .B1(_0626_),
    .A1(net527),
    .Y(_0627_),
    .A2(net483));
 sg13g2_a22oi_1 _2491_ (.Y(_0628_),
    .B1(net457),
    .B2(net12),
    .A2(net472),
    .A1(net961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2492_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0628_),
    .C1(_0503_),
    .B1(_0627_),
    .A1(_1066_),
    .Y(_0155_),
    .A2(net464));
 sg13g2_a221oi_1 _2493_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net973),
    .C1(net464),
    .B1(net483),
    .A1(net980),
    .Y(_0629_),
    .A2(net472));
 sg13g2_xnor2_1 _2494_ (.Y(_0630_),
    .A(net527),
    .B(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2495_ (.Y(_0631_),
    .B1(_0630_),
    .B2(net469),
    .A2(net457),
    .A1(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2496_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0632_),
    .VSS(VGND),
    .A1(net527),
    .A2(net460));
 sg13g2_a21oi_1 _2497_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0629_),
    .A2(_0631_),
    .Y(_0156_),
    .B1(_0632_));
 sg13g2_a221oi_1 _2498_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net967),
    .C1(net464),
    .B1(net484),
    .A1(net527),
    .Y(_0633_),
    .A2(net472));
 sg13g2_o21ai_1 _2499_ (.B1(net973),
    .VDD(VPWR),
    .Y(_0634_),
    .VSS(VGND),
    .A1(\controller.alu_buffer.buffer[6] ),
    .A2(_1285_));
 sg13g2_nand2_1 _2500_ (.Y(_0635_),
    .A(_1287_),
    .B(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2501_ (.Y(_0636_),
    .B1(_0635_),
    .B2(net468),
    .A2(net457),
    .A1(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2502_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0637_),
    .VSS(VGND),
    .A1(net973),
    .A2(net460));
 sg13g2_a21oi_1 _2503_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0633_),
    .A2(_0636_),
    .Y(_0157_),
    .B1(_0637_));
 sg13g2_a221oi_1 _2504_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.alu_buffer.buffer[10] ),
    .C1(net463),
    .B1(net483),
    .A1(\controller.alu_buffer.buffer[8] ),
    .Y(_0638_),
    .A2(net472));
 sg13g2_xnor2_1 _2505_ (.Y(_0639_),
    .A(net963),
    .B(_1288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2506_ (.Y(_0640_),
    .B1(_0639_),
    .B2(net468),
    .A2(_0607_),
    .A1(\controller.alu_buffer.buffer[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2507_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0640_),
    .C1(_0503_),
    .B1(_0638_),
    .A1(_1065_),
    .Y(_0158_),
    .A2(net463));
 sg13g2_o21ai_1 _2508_ (.B1(\controller.alu_buffer.buffer[10] ),
    .VDD(VPWR),
    .Y(_0641_),
    .VSS(VGND),
    .A1(\controller.alu_buffer.buffer[9] ),
    .A2(_1288_));
 sg13g2_nand2_1 _2509_ (.Y(_0642_),
    .A(_1290_),
    .B(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2510_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net467),
    .C1(net462),
    .B1(_0642_),
    .A1(\controller.alu_buffer.buffer[11] ),
    .Y(_0643_),
    .A2(net482));
 sg13g2_a22oi_1 _2511_ (.Y(_0644_),
    .B1(net456),
    .B2(net933),
    .A2(net471),
    .A1(\controller.alu_buffer.buffer[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2512_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0645_),
    .VSS(VGND),
    .A1(\controller.alu_buffer.buffer[10] ),
    .A2(net460));
 sg13g2_a21oi_1 _2513_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0643_),
    .A2(net934),
    .Y(_0159_),
    .B1(_0645_));
 sg13g2_a221oi_1 _2514_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net969),
    .C1(net462),
    .B1(net482),
    .A1(\controller.alu_buffer.buffer[10] ),
    .Y(_0646_),
    .A2(net471));
 sg13g2_xnor2_1 _2515_ (.Y(_0647_),
    .A(net975),
    .B(_1290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2516_ (.Y(_0648_),
    .B1(_0647_),
    .B2(net467),
    .A2(net456),
    .A1(\controller.alu_buffer.buffer[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2517_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0649_),
    .VSS(VGND),
    .A1(net975),
    .A2(net459));
 sg13g2_a21oi_1 _2518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0646_),
    .A2(_0648_),
    .Y(_0160_),
    .B1(_0649_));
 sg13g2_a221oi_1 _2519_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net954),
    .C1(net462),
    .B1(net482),
    .A1(\controller.alu_buffer.buffer[11] ),
    .Y(_0650_),
    .A2(net471));
 sg13g2_nor2_1 _2520_ (.A(\controller.alu_buffer.buffer[12] ),
    .B(_1291_),
    .Y(_0651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2521_ (.Y(_0652_),
    .A(net969),
    .B(_1291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2522_ (.Y(_0653_),
    .B1(_0652_),
    .B2(net467),
    .A2(net456),
    .A1(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2523_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0654_),
    .VSS(VGND),
    .A1(net969),
    .A2(net459));
 sg13g2_a21oi_1 _2524_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0650_),
    .A2(_0653_),
    .Y(_0161_),
    .B1(_0654_));
 sg13g2_a221oi_1 _2525_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net950),
    .C1(net462),
    .B1(net482),
    .A1(\controller.alu_buffer.buffer[12] ),
    .Y(_0655_),
    .A2(net471));
 sg13g2_nor3_1 _2526_ (.A(\controller.alu_buffer.buffer[13] ),
    .B(\controller.alu_buffer.buffer[12] ),
    .C(_1291_),
    .Y(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2527_ (.B(_0651_),
    .A(net954),
    .X(_0657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2528_ (.Y(_0658_),
    .B1(_0657_),
    .B2(net467),
    .A2(net456),
    .A1(\controller.alu_buffer.buffer[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2529_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0659_),
    .VSS(VGND),
    .A1(net954),
    .A2(net459));
 sg13g2_a21oi_1 _2530_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0655_),
    .A2(_0658_),
    .Y(_0162_),
    .B1(_0659_));
 sg13g2_nor2b_1 _2531_ (.A(_1291_),
    .B_N(_1292_),
    .Y(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2532_ (.B(_0656_),
    .A(net950),
    .X(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2533_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net466),
    .C1(net461),
    .B1(_0661_),
    .A1(net922),
    .Y(_0662_),
    .A2(net482));
 sg13g2_a22oi_1 _2534_ (.Y(_0663_),
    .B1(net455),
    .B2(net527),
    .A2(net471),
    .A1(\controller.alu_buffer.buffer[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2535_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0664_),
    .VSS(VGND),
    .A1(net950),
    .A2(net459));
 sg13g2_a21oi_1 _2536_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0662_),
    .A2(_0663_),
    .Y(_0163_),
    .B1(_0664_));
 sg13g2_a221oi_1 _2537_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.alu_buffer.buffer[16] ),
    .C1(net461),
    .B1(net481),
    .A1(\controller.alu_buffer.buffer[14] ),
    .Y(_0665_),
    .A2(net470));
 sg13g2_o21ai_1 _2538_ (.B1(_1294_),
    .VDD(VPWR),
    .Y(_0666_),
    .VSS(VGND),
    .A1(_1064_),
    .A2(_0660_));
 sg13g2_a22oi_1 _2539_ (.Y(_0667_),
    .B1(_0666_),
    .B2(net466),
    .A2(net456),
    .A1(\controller.alu_buffer.buffer[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2540_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0667_),
    .C1(_0503_),
    .B1(_0665_),
    .A1(_1064_),
    .Y(_0164_),
    .A2(net461));
 sg13g2_nor2_1 _2541_ (.A(\controller.alu_buffer.buffer[8] ),
    .B(_0562_),
    .Y(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2542_ (.A(\controller.alu_buffer.buffer[16] ),
    .B(_1294_),
    .Y(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2543_ (.A(\controller.alu_buffer.buffer[16] ),
    .B(_1294_),
    .X(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2544_ (.B1(net466),
    .VDD(VPWR),
    .Y(_0671_),
    .VSS(VGND),
    .A1(_0669_),
    .A2(_0670_));
 sg13g2_a221oi_1 _2545_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net958),
    .C1(net455),
    .B1(net481),
    .A1(net922),
    .Y(_0672_),
    .A2(net470));
 sg13g2_a21o_1 _2546_ (.A2(_0672_),
    .A1(_0671_),
    .B1(_0668_),
    .X(_0673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2547_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0674_),
    .VSS(VGND),
    .A1(net965),
    .A2(net458));
 sg13g2_a21oi_1 _2548_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net458),
    .A2(_0673_),
    .Y(_0165_),
    .B1(_0674_));
 sg13g2_a221oi_1 _2549_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net952),
    .C1(net461),
    .B1(net481),
    .A1(\controller.alu_buffer.buffer[16] ),
    .Y(_0675_),
    .A2(net470));
 sg13g2_nor3_1 _2550_ (.A(\controller.alu_buffer.buffer[17] ),
    .B(\controller.alu_buffer.buffer[16] ),
    .C(_1294_),
    .Y(_0676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2551_ (.B(_0669_),
    .A(net958),
    .X(_0677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2552_ (.Y(_0678_),
    .B1(_0677_),
    .B2(net466),
    .A2(net455),
    .A1(\controller.alu_buffer.buffer[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2553_ (.B1(net538),
    .VDD(VPWR),
    .Y(_0679_),
    .VSS(VGND),
    .A1(net958),
    .A2(net458));
 sg13g2_a21oi_1 _2554_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0675_),
    .A2(_0678_),
    .Y(_0166_),
    .B1(_0679_));
 sg13g2_nor2b_1 _2555_ (.A(\controller.alu_buffer.buffer[18] ),
    .B_N(_0676_),
    .Y(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2556_ (.B(_0676_),
    .A(net952),
    .X(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2557_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net466),
    .C1(net461),
    .B1(_0681_),
    .A1(net945),
    .Y(_0682_),
    .A2(net481));
 sg13g2_a22oi_1 _2558_ (.Y(_0683_),
    .B1(net455),
    .B2(\controller.alu_buffer.buffer[10] ),
    .A2(net470),
    .A1(\controller.alu_buffer.buffer[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2559_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0684_),
    .VSS(VGND),
    .A1(net952),
    .A2(net458));
 sg13g2_a21oi_1 _2560_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0682_),
    .A2(_0683_),
    .Y(_0167_),
    .B1(_0684_));
 sg13g2_a221oi_1 _2561_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.alu_buffer.buffer[20] ),
    .C1(net461),
    .B1(net481),
    .A1(\controller.alu_buffer.buffer[18] ),
    .Y(_0685_),
    .A2(net470));
 sg13g2_nand2b_1 _2562_ (.Y(_0686_),
    .B(net945),
    .A_N(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2563_ (.Y(_0687_),
    .B(_0686_),
    .A_N(_1296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2564_ (.Y(_0688_),
    .B1(_0687_),
    .B2(net466),
    .A2(net455),
    .A1(\controller.alu_buffer.buffer[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2565_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0689_),
    .VSS(VGND),
    .A1(net945),
    .A2(net458));
 sg13g2_a21oi_1 _2566_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0685_),
    .A2(_0688_),
    .Y(_0168_),
    .B1(_0689_));
 sg13g2_a221oi_1 _2567_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.alu_buffer.buffer[21] ),
    .C1(net461),
    .B1(net481),
    .A1(net945),
    .Y(_0690_),
    .A2(net470));
 sg13g2_xor2_1 _2568_ (.B(_1296_),
    .A(net948),
    .X(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2569_ (.Y(_0692_),
    .B1(_0691_),
    .B2(net466),
    .A2(net455),
    .A1(\controller.alu_buffer.buffer[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2570_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0693_),
    .VSS(VGND),
    .A1(net948),
    .A2(net458));
 sg13g2_a21oi_1 _2571_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0690_),
    .A2(_0692_),
    .Y(_0169_),
    .B1(_0693_));
 sg13g2_a221oi_1 _2572_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net956),
    .C1(net461),
    .B1(net481),
    .A1(net948),
    .Y(_0694_),
    .A2(net470));
 sg13g2_nor2_1 _2573_ (.A(\controller.alu_buffer.buffer[21] ),
    .B(_1297_),
    .Y(_0695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2574_ (.Y(_0696_),
    .A(net960),
    .B(_1297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2575_ (.Y(_0697_),
    .B1(_0696_),
    .B2(net466),
    .A2(net455),
    .A1(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2576_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0698_),
    .VSS(VGND),
    .A1(net960),
    .A2(net458));
 sg13g2_a21oi_1 _2577_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0694_),
    .A2(_0697_),
    .Y(_0170_),
    .B1(_0698_));
 sg13g2_nand2b_1 _2578_ (.Y(_0699_),
    .B(_0695_),
    .A_N(\controller.alu_buffer.buffer[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2579_ (.B(_0695_),
    .A(net956),
    .X(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2580_ (.Y(_0701_),
    .A(net467),
    .B(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2581_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net913),
    .C1(net456),
    .B1(net481),
    .A1(\controller.alu_buffer.buffer[21] ),
    .Y(_0702_),
    .A2(net470));
 sg13g2_nor2_1 _2582_ (.A(net950),
    .B(_0562_),
    .Y(_0703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2583_ (.A2(_0702_),
    .A1(_0701_),
    .B1(_0703_),
    .X(_0704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2584_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0705_),
    .VSS(VGND),
    .A1(net956),
    .A2(net458));
 sg13g2_a21oi_1 _2585_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net459),
    .A2(_0704_),
    .Y(_0171_),
    .B1(_0705_));
 sg13g2_a21oi_1 _2586_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net913),
    .A2(_0699_),
    .Y(_0706_),
    .B1(_1299_));
 sg13g2_nor2b_1 _2587_ (.A(_0706_),
    .B_N(net467),
    .Y(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2588_ (.A(\controller.alu_buffer.buffer[22] ),
    .B(net485),
    .C(_0561_),
    .D(_0582_),
    .X(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2589_ (.X(_0709_),
    .A(net7),
    .B(_0581_),
    .C(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2590_ (.A(net456),
    .B(_0708_),
    .C(_0709_),
    .X(_0710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2591_ (.Y(_0711_),
    .A(_1064_),
    .B(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2592_ (.B1(_0711_),
    .VDD(VPWR),
    .Y(_0712_),
    .VSS(VGND),
    .A1(_0707_),
    .A2(_0710_));
 sg13g2_o21ai_1 _2593_ (.B1(net537),
    .VDD(VPWR),
    .Y(_0713_),
    .VSS(VGND),
    .A1(net913),
    .A2(net459));
 sg13g2_a21oi_1 _2594_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net459),
    .A2(_0712_),
    .Y(_0172_),
    .B1(_0713_));
 sg13g2_and2_1 _2595_ (.A(net15),
    .B(net537),
    .X(_0173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2596_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1265_),
    .A2(_1266_),
    .Y(_0174_),
    .B1(_0503_));
 sg13g2_a21oi_1 _2597_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1267_),
    .A2(_1268_),
    .Y(_0175_),
    .B1(_0503_));
 sg13g2_o21ai_1 _2598_ (.B1(net521),
    .VDD(VPWR),
    .Y(_0714_),
    .VSS(VGND),
    .A1(_1068_),
    .A2(\controller.inst_mem.mem_data[147] ));
 sg13g2_a22oi_1 _2599_ (.Y(_0715_),
    .B1(net525),
    .B2(\controller.inst_mem.extended_word[19] ),
    .A2(net511),
    .A1(\controller.inst_mem.mem_data[171] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2600_ (.Y(_0716_),
    .B1(net496),
    .B2(\controller.inst_mem.mem_data[99] ),
    .A2(net508),
    .A1(\controller.inst_mem.mem_data[75] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2601_ (.Y(_0717_),
    .B1(net500),
    .B2(\controller.inst_mem.mem_data[123] ),
    .A2(net504),
    .A1(\controller.inst_mem.mem_data[195] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2602_ (.B(_0715_),
    .C(_0716_),
    .A(_0714_),
    .Y(_0718_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0717_));
 sg13g2_o21ai_1 _2603_ (.B1(_0718_),
    .VDD(VPWR),
    .Y(_0719_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[51] ),
    .A2(net491));
 sg13g2_or3_1 _2604_ (.A(\controller.extended_then_action[1] ),
    .B(net490),
    .C(net489),
    .X(_0720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2605_ (.B1(_0719_),
    .VDD(VPWR),
    .Y(_0721_),
    .VSS(VGND),
    .A1(net490),
    .A2(net489));
 sg13g2_and3_1 _2606_ (.X(_0722_),
    .A(net487),
    .B(_0720_),
    .C(_0721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2607_ (.Y(_0723_),
    .B1(net497),
    .B2(\controller.inst_mem.mem_data[93] ),
    .A2(net501),
    .A1(\controller.inst_mem.mem_data[117] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2608_ (.Y(_0724_),
    .B1(net526),
    .B2(\controller.extended_then_action[1] ),
    .A2(net509),
    .A1(\controller.inst_mem.mem_data[69] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2609_ (.Y(_0725_),
    .B1(_0479_),
    .B2(\controller.inst_mem.mem_data[141] ),
    .A2(net513),
    .A1(\controller.inst_mem.mem_data[165] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2610_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[189] ),
    .A2(net502),
    .Y(_0726_),
    .B1(net515));
 sg13g2_nand4_1 _2611_ (.B(_0724_),
    .C(_0725_),
    .A(_0723_),
    .Y(_0727_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0726_));
 sg13g2_o21ai_1 _2612_ (.B1(_0727_),
    .VDD(VPWR),
    .Y(_0728_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[45] ),
    .A2(net492));
 sg13g2_inv_1 _2613_ (.VDD(VPWR),
    .Y(_0729_),
    .A(_0728_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0729_),
    .Y(_0730_),
    .B1(_0485_));
 sg13g2_nor2b_1 _2615_ (.A(_0722_),
    .B_N(_0730_),
    .Y(_0731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2616_ (.Y(_0732_),
    .B(_0730_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0722_));
 sg13g2_a22oi_1 _2617_ (.Y(_0733_),
    .B1(net525),
    .B2(\controller.inst_mem.extended_word[20] ),
    .A2(net496),
    .A1(\controller.inst_mem.mem_data[100] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2618_ (.Y(_0734_),
    .B1(net508),
    .B2(\controller.inst_mem.mem_data[76] ),
    .A2(net512),
    .A1(\controller.inst_mem.mem_data[172] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2619_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[148] ),
    .C1(net518),
    .B1(net521),
    .A1(\controller.inst_mem.mem_data[124] ),
    .Y(_0735_),
    .A2(net500));
 sg13g2_nand3_1 _2620_ (.B(_0734_),
    .C(_0735_),
    .A(_0733_),
    .Y(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2621_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\controller.inst_mem.mem_data[196] ),
    .A2(net504),
    .Y(_0737_),
    .B1(_0736_));
 sg13g2_a21oi_1 _2622_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1008_),
    .A2(net518),
    .Y(_0738_),
    .B1(_0737_));
 sg13g2_mux2_1 _2623_ (.A0(\controller.extended_then_action[2] ),
    .A1(_0738_),
    .S(net488),
    .X(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2624_ (.Y(_0740_),
    .B1(net500),
    .B2(\controller.inst_mem.mem_data[118] ),
    .A2(net508),
    .A1(\controller.inst_mem.mem_data[70] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2625_ (.A2(net521),
    .A1(\controller.inst_mem.mem_data[142] ),
    .B1(_1231_),
    .X(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2626_ (.Y(_0742_),
    .B1(net496),
    .B2(\controller.inst_mem.mem_data[94] ),
    .A2(net512),
    .A1(\controller.inst_mem.mem_data[166] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2627_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.extended_then_action[2] ),
    .C1(_0741_),
    .B1(net525),
    .A1(\controller.inst_mem.mem_data[190] ),
    .Y(_0743_),
    .A2(net504));
 sg13g2_nand3_1 _2628_ (.B(_0742_),
    .C(_0743_),
    .A(_0740_),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2629_ (.B1(_0744_),
    .VDD(VPWR),
    .Y(_0745_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[46] ),
    .A2(net492));
 sg13g2_o21ai_1 _2630_ (.B1(_0486_),
    .VDD(VPWR),
    .Y(_0746_),
    .VSS(VGND),
    .A1(net487),
    .A2(_0745_));
 sg13g2_a21oi_2 _2631_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0746_),
    .Y(_0747_),
    .A2(_0739_),
    .A1(net487));
 sg13g2_a21o_2 _2632_ (.A2(_0739_),
    .A1(net487),
    .B1(_0746_),
    .X(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2633_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[146] ),
    .C1(net518),
    .B1(net521),
    .A1(\controller.inst_mem.mem_data[170] ),
    .Y(_0749_),
    .A2(net512));
 sg13g2_a22oi_1 _2634_ (.Y(_0750_),
    .B1(net500),
    .B2(\controller.inst_mem.mem_data[122] ),
    .A2(net504),
    .A1(\controller.inst_mem.mem_data[194] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2635_ (.Y(_0751_),
    .B1(net525),
    .B2(\controller.inst_mem.extended_word[18] ),
    .A2(net496),
    .A1(\controller.inst_mem.mem_data[98] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2636_ (.B(_0750_),
    .C(_0751_),
    .A(_0749_),
    .Y(_0752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2637_ (.A2(net508),
    .A1(\controller.inst_mem.mem_data[74] ),
    .B1(_0752_),
    .X(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2638_ (.B1(_0753_),
    .VDD(VPWR),
    .Y(_0754_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[50] ),
    .A2(net491));
 sg13g2_o21ai_1 _2639_ (.B1(_0754_),
    .VDD(VPWR),
    .Y(_0755_),
    .VSS(VGND),
    .A1(net490),
    .A2(net489));
 sg13g2_or3_1 _2640_ (.A(\controller.extended_then_action[0] ),
    .B(net490),
    .C(net489),
    .X(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2641_ (.B(_0755_),
    .C(_0756_),
    .A(net487),
    .Y(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2642_ (.Y(_0758_),
    .A(_1016_),
    .B(net516),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2643_ (.A2(net519),
    .A1(\controller.inst_mem.mem_data[140] ),
    .B1(net515),
    .X(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2644_ (.Y(_0760_),
    .B1(net526),
    .B2(\controller.extended_then_action[0] ),
    .A2(net505),
    .A1(\controller.inst_mem.mem_data[188] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2645_ (.Y(_0761_),
    .B1(net494),
    .B2(\controller.inst_mem.mem_data[92] ),
    .A2(net509),
    .A1(\controller.inst_mem.mem_data[68] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2646_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\controller.inst_mem.mem_data[116] ),
    .C1(_0759_),
    .B1(net501),
    .A1(\controller.inst_mem.mem_data[164] ),
    .Y(_0762_),
    .A2(net513));
 sg13g2_nand3_1 _2647_ (.B(_0761_),
    .C(_0762_),
    .A(_0760_),
    .Y(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2648_ (.B(_0758_),
    .C(_0763_),
    .A(_0475_),
    .Y(_0764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2649_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0485_),
    .Y(_0765_),
    .A2(_0764_),
    .A1(_0757_));
 sg13g2_nor2_1 _2650_ (.A(_0747_),
    .B(_0765_),
    .Y(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2651_ (.B1(_0732_),
    .VDD(VPWR),
    .Y(_0767_),
    .VSS(VGND),
    .A1(_0747_),
    .A2(_0765_));
 sg13g2_and2_1 _2652_ (.A(_0747_),
    .B(_0765_),
    .X(_0768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2653_ (.Y(_0769_),
    .A(net474),
    .B(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2654_ (.A(_0767_),
    .B(_0768_),
    .Y(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2655_ (.Y(_0771_),
    .B(net448),
    .A_N(net947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2656_ (.A0(_0766_),
    .A1(_0769_),
    .S(net480),
    .X(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2657_ (.B1(_0767_),
    .VDD(VPWR),
    .Y(_0773_),
    .VSS(VGND),
    .A1(_0732_),
    .A2(_0769_));
 sg13g2_and2_1 _2658_ (.A(_0732_),
    .B(_0768_),
    .X(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2659_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net7),
    .C1(net447),
    .B1(_0774_),
    .A1(net671),
    .Y(_0775_),
    .A2(net479));
 sg13g2_o21ai_1 _2660_ (.B1(net540),
    .VDD(VPWR),
    .Y(_0776_),
    .VSS(VGND),
    .A1(net947),
    .A2(net444));
 sg13g2_a21oi_1 _2661_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0771_),
    .A2(_0775_),
    .Y(_0176_),
    .B1(_0776_));
 sg13g2_and2_1 _2662_ (.A(net930),
    .B(\controller.counter2.counter_0[0] ),
    .X(_0777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2663_ (.B1(net448),
    .VDD(VPWR),
    .Y(_0778_),
    .VSS(VGND),
    .A1(_0405_),
    .A2(_0777_));
 sg13g2_a221oi_1 _2664_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net8),
    .C1(net446),
    .B1(_0774_),
    .A1(net695),
    .Y(_0779_),
    .A2(net479));
 sg13g2_o21ai_1 _2665_ (.B1(net540),
    .VDD(VPWR),
    .Y(_0780_),
    .VSS(VGND),
    .A1(net930),
    .A2(net444));
 sg13g2_a21oi_1 _2666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0778_),
    .A2(_0779_),
    .Y(_0177_),
    .B1(_0780_));
 sg13g2_nor2b_1 _2667_ (.A(_0405_),
    .B_N(net919),
    .Y(_0781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2668_ (.B1(net448),
    .VDD(VPWR),
    .Y(_0782_),
    .VSS(VGND),
    .A1(_0406_),
    .A2(_0781_));
 sg13g2_a221oi_1 _2669_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net9),
    .C1(net446),
    .B1(_0774_),
    .A1(net832),
    .Y(_0783_),
    .A2(net479));
 sg13g2_o21ai_1 _2670_ (.B1(net540),
    .VDD(VPWR),
    .Y(_0784_),
    .VSS(VGND),
    .A1(net919),
    .A2(net444));
 sg13g2_a21oi_1 _2671_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0782_),
    .A2(_0783_),
    .Y(_0178_),
    .B1(_0784_));
 sg13g2_xnor2_1 _2672_ (.Y(_0785_),
    .A(net928),
    .B(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2673_ (.Y(_0786_),
    .B(net448),
    .A_N(_0785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2674_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net10),
    .C1(net446),
    .B1(_0774_),
    .A1(net838),
    .Y(_0787_),
    .A2(net479));
 sg13g2_o21ai_1 _2675_ (.B1(net540),
    .VDD(VPWR),
    .Y(_0788_),
    .VSS(VGND),
    .A1(net928),
    .A2(net444));
 sg13g2_a21oi_1 _2676_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0786_),
    .A2(_0787_),
    .Y(_0179_),
    .B1(_0788_));
 sg13g2_and2_1 _2677_ (.A(net944),
    .B(_0407_),
    .X(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2678_ (.B1(net448),
    .VDD(VPWR),
    .Y(_0790_),
    .VSS(VGND),
    .A1(_0408_),
    .A2(_0789_));
 sg13g2_a221oi_1 _2679_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net11),
    .C1(net446),
    .B1(_0774_),
    .A1(net419),
    .Y(_0791_),
    .A2(net479));
 sg13g2_o21ai_1 _2680_ (.B1(net540),
    .VDD(VPWR),
    .Y(_0792_),
    .VSS(VGND),
    .A1(net944),
    .A2(net444));
 sg13g2_a21oi_1 _2681_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0790_),
    .A2(_0791_),
    .Y(_0180_),
    .B1(_0792_));
 sg13g2_nor2b_1 _2682_ (.A(_0408_),
    .B_N(net938),
    .Y(_0793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2683_ (.B1(net448),
    .VDD(VPWR),
    .Y(_0794_),
    .VSS(VGND),
    .A1(_0409_),
    .A2(_0793_));
 sg13g2_a221oi_1 _2684_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net12),
    .C1(net446),
    .B1(_0774_),
    .A1(net774),
    .Y(_0795_),
    .A2(net479));
 sg13g2_o21ai_1 _2685_ (.B1(net540),
    .VDD(VPWR),
    .Y(_0796_),
    .VSS(VGND),
    .A1(net938),
    .A2(net444));
 sg13g2_a21oi_1 _2686_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0794_),
    .A2(_0795_),
    .Y(_0181_),
    .B1(_0796_));
 sg13g2_nor2b_1 _2687_ (.A(_0409_),
    .B_N(net894),
    .Y(_0797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2688_ (.B1(net448),
    .VDD(VPWR),
    .Y(_0798_),
    .VSS(VGND),
    .A1(_0410_),
    .A2(_0797_));
 sg13g2_a221oi_1 _2689_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net13),
    .C1(net446),
    .B1(_0774_),
    .A1(net715),
    .Y(_0799_),
    .A2(net479));
 sg13g2_o21ai_1 _2690_ (.B1(net539),
    .VDD(VPWR),
    .Y(_0800_),
    .VSS(VGND),
    .A1(net894),
    .A2(net444));
 sg13g2_a21oi_1 _2691_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0798_),
    .A2(_0799_),
    .Y(_0182_),
    .B1(_0800_));
 sg13g2_xnor2_1 _2692_ (.Y(_0801_),
    .A(_1063_),
    .B(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2693_ (.Y(_0802_),
    .A(net449),
    .B(_0801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2694_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net14),
    .C1(net446),
    .B1(_0774_),
    .A1(net824),
    .Y(_0803_),
    .A2(net479));
 sg13g2_a221oi_1 _2695_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0803_),
    .C1(_0503_),
    .B1(_0802_),
    .A1(_1063_),
    .Y(_0183_),
    .A2(net447));
 sg13g2_xnor2_1 _2696_ (.Y(_0804_),
    .A(net896),
    .B(_0411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2697_ (.Y(_0805_),
    .B1(net448),
    .B2(_0804_),
    .A2(_0767_),
    .A1(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2698_ (.B1(net541),
    .VDD(VPWR),
    .Y(_0806_),
    .VSS(VGND),
    .A1(net896),
    .A2(net444));
 sg13g2_a21oi_1 _2699_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net445),
    .A2(_0805_),
    .Y(_0184_),
    .B1(_0806_));
 sg13g2_o21ai_1 _2700_ (.B1(net886),
    .VDD(VPWR),
    .Y(_0807_),
    .VSS(VGND),
    .A1(\controller.counter2.counter_0[8] ),
    .A2(_0411_));
 sg13g2_nand2_1 _2701_ (.Y(_0808_),
    .A(_0413_),
    .B(_0807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2702_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0808_),
    .C1(net446),
    .B1(net449),
    .A1(net390),
    .Y(_0809_),
    .A2(net480));
 sg13g2_o21ai_1 _2703_ (.B1(net541),
    .VDD(VPWR),
    .Y(_0810_),
    .VSS(VGND),
    .A1(net886),
    .A2(net445));
 sg13g2_nor2_1 _2704_ (.A(_0809_),
    .B(_0810_),
    .Y(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2705_ (.Y(_0811_),
    .A(net924),
    .B(_0413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2706_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0811_),
    .C1(net447),
    .B1(net449),
    .A1(net713),
    .Y(_0812_),
    .A2(net480));
 sg13g2_o21ai_1 _2707_ (.B1(net541),
    .VDD(VPWR),
    .Y(_0813_),
    .VSS(VGND),
    .A1(net924),
    .A2(_0773_));
 sg13g2_nor2_1 _2708_ (.A(_0812_),
    .B(_0813_),
    .Y(_0186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2709_ (.Y(_0814_),
    .A(net897),
    .B(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2710_ (.Y(_0815_),
    .B1(net449),
    .B2(_0814_),
    .A2(_0767_),
    .A1(net681),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2711_ (.B1(net541),
    .VDD(VPWR),
    .Y(_0816_),
    .VSS(VGND),
    .A1(net897),
    .A2(net445));
 sg13g2_a21oi_1 _2712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net445),
    .A2(_0815_),
    .Y(_0187_),
    .B1(_0816_));
 sg13g2_xnor2_1 _2713_ (.Y(_0817_),
    .A(net916),
    .B(_0415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2714_ (.Y(_0818_),
    .B1(net449),
    .B2(_0817_),
    .A2(_0767_),
    .A1(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2715_ (.B1(net541),
    .VDD(VPWR),
    .Y(_0819_),
    .VSS(VGND),
    .A1(net916),
    .A2(net445));
 sg13g2_a21oi_1 _2716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net445),
    .A2(_0818_),
    .Y(_0188_),
    .B1(_0819_));
 sg13g2_o21ai_1 _2717_ (.B1(net899),
    .VDD(VPWR),
    .Y(_0820_),
    .VSS(VGND),
    .A1(\controller.counter2.counter_0[12] ),
    .A2(_0415_));
 sg13g2_nand2b_1 _2718_ (.Y(_0821_),
    .B(_0820_),
    .A_N(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2719_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0821_),
    .C1(net447),
    .B1(net449),
    .A1(net707),
    .Y(_0822_),
    .A2(net480));
 sg13g2_o21ai_1 _2720_ (.B1(net542),
    .VDD(VPWR),
    .Y(_0823_),
    .VSS(VGND),
    .A1(net899),
    .A2(_0773_));
 sg13g2_nor2_1 _2721_ (.A(_0822_),
    .B(_0823_),
    .Y(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2722_ (.B(_0417_),
    .A(net893),
    .X(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2723_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0824_),
    .C1(net447),
    .B1(net449),
    .A1(net694),
    .Y(_0825_),
    .A2(net480));
 sg13g2_o21ai_1 _2724_ (.B1(net542),
    .VDD(VPWR),
    .Y(_0826_),
    .VSS(VGND),
    .A1(net893),
    .A2(_0773_));
 sg13g2_nor2_1 _2725_ (.A(_0825_),
    .B(_0826_),
    .Y(_0190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2726_ (.B(_0418_),
    .A(net906),
    .X(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2727_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0827_),
    .C1(net447),
    .B1(_0770_),
    .A1(net348),
    .Y(_0828_),
    .A2(net480));
 sg13g2_o21ai_1 _2728_ (.B1(net541),
    .VDD(VPWR),
    .Y(_0829_),
    .VSS(VGND),
    .A1(net906),
    .A2(net445));
 sg13g2_nor2_1 _2729_ (.A(_0828_),
    .B(_0829_),
    .Y(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2730_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0830_),
    .B(_0765_),
    .A(net480));
 sg13g2_nor2_1 _2731_ (.A(net892),
    .B(net451),
    .Y(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2732_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net418),
    .A2(net451),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_o21ai_1 _2733_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0833_),
    .VSS(VGND),
    .A1(net892),
    .A2(net475));
 sg13g2_a21oi_1 _2734_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net475),
    .A2(_0832_),
    .Y(_0192_),
    .B1(_0833_));
 sg13g2_xor2_1 _2735_ (.B(net892),
    .A(net915),
    .X(_0834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2736_ (.A(net454),
    .B(_0834_),
    .Y(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2737_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net410),
    .A2(net454),
    .Y(_0836_),
    .B1(_0835_));
 sg13g2_o21ai_1 _2738_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0837_),
    .VSS(VGND),
    .A1(net915),
    .A2(net475));
 sg13g2_a21oi_1 _2739_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net475),
    .A2(_0836_),
    .Y(_0193_),
    .B1(_0837_));
 sg13g2_o21ai_1 _2740_ (.B1(net911),
    .VDD(VPWR),
    .Y(_0838_),
    .VSS(VGND),
    .A1(\controller.counter2.counter_1[1] ),
    .A2(\controller.counter2.counter_1[0] ));
 sg13g2_nor2b_1 _2741_ (.A(_1269_),
    .B_N(_0838_),
    .Y(_0839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2742_ (.A(net454),
    .B(_0839_),
    .Y(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2743_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net409),
    .A2(net451),
    .Y(_0841_),
    .B1(_0840_));
 sg13g2_o21ai_1 _2744_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0842_),
    .VSS(VGND),
    .A1(net911),
    .A2(net475));
 sg13g2_a21oi_1 _2745_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net475),
    .A2(_0841_),
    .Y(_0194_),
    .B1(_0842_));
 sg13g2_nand2b_1 _2746_ (.Y(_0843_),
    .B(net890),
    .A_N(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2747_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1270_),
    .A2(_0843_),
    .Y(_0844_),
    .B1(net451));
 sg13g2_a21oi_1 _2748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net344),
    .A2(net451),
    .Y(_0845_),
    .B1(_0844_));
 sg13g2_o21ai_1 _2749_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0846_),
    .VSS(VGND),
    .A1(net890),
    .A2(net477));
 sg13g2_a21oi_1 _2750_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net477),
    .A2(_0845_),
    .Y(_0195_),
    .B1(_0846_));
 sg13g2_xor2_1 _2751_ (.B(_1270_),
    .A(net903),
    .X(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2752_ (.A(net452),
    .B(_0847_),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net736),
    .A2(net452),
    .Y(_0849_),
    .B1(_0848_));
 sg13g2_o21ai_1 _2754_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0850_),
    .VSS(VGND),
    .A1(net903),
    .A2(net476));
 sg13g2_a21oi_1 _2755_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net476),
    .A2(_0849_),
    .Y(_0196_),
    .B1(_0850_));
 sg13g2_o21ai_1 _2756_ (.B1(net910),
    .VDD(VPWR),
    .Y(_0851_),
    .VSS(VGND),
    .A1(net903),
    .A2(_1270_));
 sg13g2_a21oi_1 _2757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1271_),
    .A2(_0851_),
    .Y(_0852_),
    .B1(net452));
 sg13g2_a21oi_1 _2758_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net718),
    .A2(net453),
    .Y(_0853_),
    .B1(_0852_));
 sg13g2_o21ai_1 _2759_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(net910),
    .A2(net476));
 sg13g2_a21oi_1 _2760_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net476),
    .A2(_0853_),
    .Y(_0197_),
    .B1(_0854_));
 sg13g2_nand2_1 _2761_ (.Y(_0855_),
    .A(net888),
    .B(_1271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2762_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1272_),
    .A2(_0855_),
    .Y(_0856_),
    .B1(net452));
 sg13g2_a21oi_1 _2763_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net840),
    .A2(net453),
    .Y(_0857_),
    .B1(_0856_));
 sg13g2_o21ai_1 _2764_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0858_),
    .VSS(VGND),
    .A1(net888),
    .A2(net477));
 sg13g2_a21oi_1 _2765_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net477),
    .A2(_0857_),
    .Y(_0198_),
    .B1(_0858_));
 sg13g2_nand2_1 _2766_ (.Y(_0859_),
    .A(net932),
    .B(_1272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2767_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1273_),
    .A2(_0859_),
    .Y(_0860_),
    .B1(net452));
 sg13g2_a21oi_1 _2768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net820),
    .A2(net452),
    .Y(_0861_),
    .B1(_0860_));
 sg13g2_o21ai_1 _2769_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0862_),
    .VSS(VGND),
    .A1(net932),
    .A2(net476));
 sg13g2_a21oi_1 _2770_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net476),
    .A2(_0861_),
    .Y(_0199_),
    .B1(_0862_));
 sg13g2_xor2_1 _2771_ (.B(_1273_),
    .A(net921),
    .X(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2772_ (.A(net452),
    .B(_0863_),
    .Y(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net811),
    .A2(net452),
    .Y(_0865_),
    .B1(_0864_));
 sg13g2_o21ai_1 _2774_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0866_),
    .VSS(VGND),
    .A1(net921),
    .A2(net476));
 sg13g2_a21oi_1 _2775_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net476),
    .A2(_0865_),
    .Y(_0200_),
    .B1(_0866_));
 sg13g2_o21ai_1 _2776_ (.B1(net901),
    .VDD(VPWR),
    .Y(_0867_),
    .VSS(VGND),
    .A1(\controller.counter2.counter_1[8] ),
    .A2(_1273_));
 sg13g2_nor2b_1 _2777_ (.A(_1274_),
    .B_N(_0867_),
    .Y(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2778_ (.A(net453),
    .B(_0868_),
    .Y(_0869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2779_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net687),
    .A2(net453),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_o21ai_1 _2780_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0871_),
    .VSS(VGND),
    .A1(net901),
    .A2(net478));
 sg13g2_a21oi_1 _2781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net478),
    .A2(_0870_),
    .Y(_0201_),
    .B1(_0871_));
 sg13g2_nand2b_1 _2782_ (.Y(_0872_),
    .B(net907),
    .A_N(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2783_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1275_),
    .A2(_0872_),
    .Y(_0873_),
    .B1(net453));
 sg13g2_a21oi_1 _2784_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net818),
    .A2(net453),
    .Y(_0874_),
    .B1(_0873_));
 sg13g2_o21ai_1 _2785_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0875_),
    .VSS(VGND),
    .A1(net907),
    .A2(net478));
 sg13g2_a21oi_1 _2786_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net478),
    .A2(_0874_),
    .Y(_0202_),
    .B1(_0875_));
 sg13g2_nand2_1 _2787_ (.Y(_0876_),
    .A(net883),
    .B(_1275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2788_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1277_),
    .A2(_0876_),
    .Y(_0877_),
    .B1(net451));
 sg13g2_a21oi_1 _2789_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net396),
    .A2(net451),
    .Y(_0878_),
    .B1(_0877_));
 sg13g2_o21ai_1 _2790_ (.B1(net543),
    .VDD(VPWR),
    .Y(_0879_),
    .VSS(VGND),
    .A1(net883),
    .A2(net478));
 sg13g2_a21oi_1 _2791_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net478),
    .A2(_0878_),
    .Y(_0203_),
    .B1(_0879_));
 sg13g2_xor2_1 _2792_ (.B(_1277_),
    .A(net942),
    .X(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2793_ (.A(net450),
    .B(_0880_),
    .Y(_0881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2794_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net822),
    .A2(net450),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_o21ai_1 _2795_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0883_),
    .VSS(VGND),
    .A1(net942),
    .A2(net474));
 sg13g2_a21oi_1 _2796_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net474),
    .A2(_0882_),
    .Y(_0204_),
    .B1(_0883_));
 sg13g2_nor3_1 _2797_ (.A(net926),
    .B(\controller.counter2.counter_1[12] ),
    .C(_1277_),
    .Y(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2798_ (.B1(net926),
    .VDD(VPWR),
    .Y(_0885_),
    .VSS(VGND),
    .A1(\controller.counter2.counter_1[12] ),
    .A2(_1277_));
 sg13g2_nor2b_1 _2799_ (.A(_0884_),
    .B_N(_0885_),
    .Y(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2800_ (.A(net450),
    .B(_0886_),
    .Y(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2801_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net440),
    .A2(net450),
    .Y(_0888_),
    .B1(_0887_));
 sg13g2_o21ai_1 _2802_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0889_),
    .VSS(VGND),
    .A1(net926),
    .A2(net474));
 sg13g2_a21oi_1 _2803_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net475),
    .A2(_0888_),
    .Y(_0205_),
    .B1(_0889_));
 sg13g2_nand2b_1 _2804_ (.Y(_0890_),
    .B(_0884_),
    .A_N(net904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2805_ (.Y(_0891_),
    .A(net904),
    .B(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2806_ (.A(net450),
    .B(_0891_),
    .Y(_0892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2807_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net689),
    .A2(net450),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_o21ai_1 _2808_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0894_),
    .VSS(VGND),
    .A1(net904),
    .A2(net474));
 sg13g2_a21oi_1 _2809_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net474),
    .A2(_0893_),
    .Y(_0206_),
    .B1(_0894_));
 sg13g2_a21oi_1 _2810_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net909),
    .A2(_0890_),
    .Y(_0895_),
    .B1(_1279_));
 sg13g2_nor2_1 _2811_ (.A(net450),
    .B(_0895_),
    .Y(_0896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2812_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net873),
    .A2(net450),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_o21ai_1 _2813_ (.B1(net544),
    .VDD(VPWR),
    .Y(_0898_),
    .VSS(VGND),
    .A1(net909),
    .A2(net474));
 sg13g2_a21oi_1 _2814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net474),
    .A2(_0897_),
    .Y(_0207_),
    .B1(_0898_));
 sg13g2_o21ai_1 _2815_ (.B1(net637),
    .VDD(VPWR),
    .Y(_0899_),
    .VSS(VGND),
    .A1(net671),
    .A2(net580));
 sg13g2_a21oi_1 _2816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1061_),
    .A2(net580),
    .Y(_0208_),
    .B1(_0899_));
 sg13g2_o21ai_1 _2817_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0900_),
    .VSS(VGND),
    .A1(\controller.const_data[1] ),
    .A2(net570));
 sg13g2_a21oi_1 _2818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1060_),
    .A2(net570),
    .Y(_0209_),
    .B1(_0900_));
 sg13g2_o21ai_1 _2819_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0901_),
    .VSS(VGND),
    .A1(\controller.const_data[2] ),
    .A2(net570));
 sg13g2_a21oi_1 _2820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1059_),
    .A2(net570),
    .Y(_0210_),
    .B1(_0901_));
 sg13g2_o21ai_1 _2821_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0902_),
    .VSS(VGND),
    .A1(\controller.const_data[3] ),
    .A2(net570));
 sg13g2_a21oi_1 _2822_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1058_),
    .A2(net570),
    .Y(_0211_),
    .B1(_0902_));
 sg13g2_o21ai_1 _2823_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0903_),
    .VSS(VGND),
    .A1(net419),
    .A2(net569));
 sg13g2_a21oi_1 _2824_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1057_),
    .A2(net569),
    .Y(_0212_),
    .B1(_0903_));
 sg13g2_o21ai_1 _2825_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0904_),
    .VSS(VGND),
    .A1(\controller.const_data[5] ),
    .A2(net569));
 sg13g2_a21oi_1 _2826_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1056_),
    .A2(net569),
    .Y(_0213_),
    .B1(_0904_));
 sg13g2_o21ai_1 _2827_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0905_),
    .VSS(VGND),
    .A1(net715),
    .A2(net569));
 sg13g2_a21oi_1 _2828_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1055_),
    .A2(net569),
    .Y(_0214_),
    .B1(_0905_));
 sg13g2_o21ai_1 _2829_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0906_),
    .VSS(VGND),
    .A1(\controller.const_data[7] ),
    .A2(net569));
 sg13g2_a21oi_1 _2830_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1054_),
    .A2(net569),
    .Y(_0215_),
    .B1(_0906_));
 sg13g2_o21ai_1 _2831_ (.B1(net637),
    .VDD(VPWR),
    .Y(_0907_),
    .VSS(VGND),
    .A1(net788),
    .A2(net571));
 sg13g2_a21oi_1 _2832_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1053_),
    .A2(net570),
    .Y(_0216_),
    .B1(_0907_));
 sg13g2_o21ai_1 _2833_ (.B1(net637),
    .VDD(VPWR),
    .Y(_0908_),
    .VSS(VGND),
    .A1(net390),
    .A2(net571));
 sg13g2_a21oi_1 _2834_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1052_),
    .A2(net571),
    .Y(_0217_),
    .B1(_0908_));
 sg13g2_o21ai_1 _2835_ (.B1(net636),
    .VDD(VPWR),
    .Y(_0909_),
    .VSS(VGND),
    .A1(\controller.const_data[10] ),
    .A2(net571));
 sg13g2_a21oi_1 _2836_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1051_),
    .A2(net571),
    .Y(_0218_),
    .B1(_0909_));
 sg13g2_o21ai_1 _2837_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0910_),
    .VSS(VGND),
    .A1(net681),
    .A2(net571));
 sg13g2_a21oi_1 _2838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1050_),
    .A2(net571),
    .Y(_0219_),
    .B1(_0910_));
 sg13g2_o21ai_1 _2839_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0911_),
    .VSS(VGND),
    .A1(net372),
    .A2(net577));
 sg13g2_a21oi_1 _2840_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1049_),
    .A2(net577),
    .Y(_0220_),
    .B1(_0911_));
 sg13g2_o21ai_1 _2841_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0912_),
    .VSS(VGND),
    .A1(\controller.const_data[13] ),
    .A2(net577));
 sg13g2_a21oi_1 _2842_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1048_),
    .A2(net577),
    .Y(_0221_),
    .B1(_0912_));
 sg13g2_o21ai_1 _2843_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0913_),
    .VSS(VGND),
    .A1(net694),
    .A2(net577));
 sg13g2_a21oi_1 _2844_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1047_),
    .A2(net577),
    .Y(_0222_),
    .B1(_0913_));
 sg13g2_o21ai_1 _2845_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0914_),
    .VSS(VGND),
    .A1(net348),
    .A2(net577));
 sg13g2_a21oi_1 _2846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1046_),
    .A2(net577),
    .Y(_0223_),
    .B1(_0914_));
 sg13g2_o21ai_1 _2847_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0915_),
    .VSS(VGND),
    .A1(\controller.const_data[16] ),
    .A2(net578));
 sg13g2_a21oi_1 _2848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1045_),
    .A2(net578),
    .Y(_0224_),
    .B1(_0915_));
 sg13g2_o21ai_1 _2849_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0916_),
    .VSS(VGND),
    .A1(net410),
    .A2(net576));
 sg13g2_a21oi_1 _2850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1044_),
    .A2(net576),
    .Y(_0225_),
    .B1(_0916_));
 sg13g2_o21ai_1 _2851_ (.B1(net640),
    .VDD(VPWR),
    .Y(_0917_),
    .VSS(VGND),
    .A1(net409),
    .A2(net576));
 sg13g2_a21oi_1 _2852_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1043_),
    .A2(net578),
    .Y(_0226_),
    .B1(_0917_));
 sg13g2_o21ai_1 _2853_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0918_),
    .VSS(VGND),
    .A1(net344),
    .A2(net612));
 sg13g2_a21oi_1 _2854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1042_),
    .A2(net576),
    .Y(_0227_),
    .B1(_0918_));
 sg13g2_o21ai_1 _2855_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0919_),
    .VSS(VGND),
    .A1(\controller.const_data[20] ),
    .A2(net612));
 sg13g2_a21oi_1 _2856_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1041_),
    .A2(net612),
    .Y(_0228_),
    .B1(_0919_));
 sg13g2_o21ai_1 _2857_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0920_),
    .VSS(VGND),
    .A1(net718),
    .A2(net612));
 sg13g2_a21oi_1 _2858_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1040_),
    .A2(net614),
    .Y(_0229_),
    .B1(_0920_));
 sg13g2_o21ai_1 _2859_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(\controller.const_data[22] ),
    .A2(net613));
 sg13g2_a21oi_1 _2860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1039_),
    .A2(net613),
    .Y(_0230_),
    .B1(_0921_));
 sg13g2_o21ai_1 _2861_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0922_),
    .VSS(VGND),
    .A1(net820),
    .A2(net614));
 sg13g2_a21oi_1 _2862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1038_),
    .A2(net613),
    .Y(_0231_),
    .B1(_0922_));
 sg13g2_o21ai_1 _2863_ (.B1(net659),
    .VDD(VPWR),
    .Y(_0923_),
    .VSS(VGND),
    .A1(net811),
    .A2(net613));
 sg13g2_a21oi_1 _2864_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1037_),
    .A2(net614),
    .Y(_0232_),
    .B1(_0923_));
 sg13g2_o21ai_1 _2865_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0924_),
    .VSS(VGND),
    .A1(net687),
    .A2(net613));
 sg13g2_a21oi_1 _2866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1036_),
    .A2(net613),
    .Y(_0233_),
    .B1(_0924_));
 sg13g2_o21ai_1 _2867_ (.B1(net659),
    .VDD(VPWR),
    .Y(_0925_),
    .VSS(VGND),
    .A1(\controller.const_data[26] ),
    .A2(net613));
 sg13g2_a21oi_1 _2868_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1035_),
    .A2(net613),
    .Y(_0234_),
    .B1(_0925_));
 sg13g2_o21ai_1 _2869_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0926_),
    .VSS(VGND),
    .A1(net396),
    .A2(net612));
 sg13g2_a21oi_1 _2870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1034_),
    .A2(net612),
    .Y(_0235_),
    .B1(_0926_));
 sg13g2_o21ai_1 _2871_ (.B1(net658),
    .VDD(VPWR),
    .Y(_0927_),
    .VSS(VGND),
    .A1(\controller.const_data[28] ),
    .A2(net612));
 sg13g2_a21oi_1 _2872_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1033_),
    .A2(net612),
    .Y(_0236_),
    .B1(_0927_));
 sg13g2_o21ai_1 _2873_ (.B1(net641),
    .VDD(VPWR),
    .Y(_0928_),
    .VSS(VGND),
    .A1(net440),
    .A2(net576));
 sg13g2_a21oi_1 _2874_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1032_),
    .A2(net576),
    .Y(_0237_),
    .B1(_0928_));
 sg13g2_o21ai_1 _2875_ (.B1(net641),
    .VDD(VPWR),
    .Y(_0929_),
    .VSS(VGND),
    .A1(\controller.const_data[30] ),
    .A2(net576));
 sg13g2_a21oi_1 _2876_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1031_),
    .A2(net576),
    .Y(_0238_),
    .B1(_0929_));
 sg13g2_o21ai_1 _2877_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0930_),
    .VSS(VGND),
    .A1(\controller.const_data[31] ),
    .A2(net574));
 sg13g2_a21oi_1 _2878_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1030_),
    .A2(net574),
    .Y(_0239_),
    .B1(_0930_));
 sg13g2_o21ai_1 _2879_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0931_),
    .VSS(VGND),
    .A1(net777),
    .A2(net590));
 sg13g2_a21oi_1 _2880_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1029_),
    .A2(net590),
    .Y(_0240_),
    .B1(_0931_));
 sg13g2_o21ai_1 _2881_ (.B1(net644),
    .VDD(VPWR),
    .Y(_0932_),
    .VSS(VGND),
    .A1(net720),
    .A2(net587));
 sg13g2_a21oi_1 _2882_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1028_),
    .A2(net587),
    .Y(_0241_),
    .B1(_0932_));
 sg13g2_o21ai_1 _2883_ (.B1(net642),
    .VDD(VPWR),
    .Y(_0933_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[34] ),
    .A2(net582));
 sg13g2_a21oi_1 _2884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1027_),
    .A2(net583),
    .Y(_0242_),
    .B1(_0933_));
 sg13g2_o21ai_1 _2885_ (.B1(net642),
    .VDD(VPWR),
    .Y(_0934_),
    .VSS(VGND),
    .A1(net748),
    .A2(net582));
 sg13g2_a21oi_1 _2886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1026_),
    .A2(net582),
    .Y(_0243_),
    .B1(_0934_));
 sg13g2_o21ai_1 _2887_ (.B1(net645),
    .VDD(VPWR),
    .Y(_0935_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[36] ),
    .A2(net561));
 sg13g2_a21oi_1 _2888_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1025_),
    .A2(net582),
    .Y(_0244_),
    .B1(_0935_));
 sg13g2_o21ai_1 _2889_ (.B1(net631),
    .VDD(VPWR),
    .Y(_0936_),
    .VSS(VGND),
    .A1(net869),
    .A2(net561));
 sg13g2_a21oi_1 _2890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1024_),
    .A2(net561),
    .Y(_0245_),
    .B1(_0936_));
 sg13g2_o21ai_1 _2891_ (.B1(net631),
    .VDD(VPWR),
    .Y(_0937_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[38] ),
    .A2(net558));
 sg13g2_a21oi_1 _2892_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1023_),
    .A2(net558),
    .Y(_0246_),
    .B1(_0937_));
 sg13g2_o21ai_1 _2893_ (.B1(net626),
    .VDD(VPWR),
    .Y(_0938_),
    .VSS(VGND),
    .A1(net799),
    .A2(net547));
 sg13g2_a21oi_1 _2894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1022_),
    .A2(net551),
    .Y(_0247_),
    .B1(_0938_));
 sg13g2_o21ai_1 _2895_ (.B1(net627),
    .VDD(VPWR),
    .Y(_0939_),
    .VSS(VGND),
    .A1(net722),
    .A2(net547));
 sg13g2_a21oi_1 _2896_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1021_),
    .A2(net547),
    .Y(_0248_),
    .B1(_0939_));
 sg13g2_o21ai_1 _2897_ (.B1(net635),
    .VDD(VPWR),
    .Y(_0940_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[41] ),
    .A2(net554));
 sg13g2_a21oi_1 _2898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1020_),
    .A2(net554),
    .Y(_0249_),
    .B1(_0940_));
 sg13g2_o21ai_1 _2899_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0941_),
    .VSS(VGND),
    .A1(net740),
    .A2(net563));
 sg13g2_a21oi_1 _2900_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1019_),
    .A2(net563),
    .Y(_0250_),
    .B1(_0941_));
 sg13g2_o21ai_1 _2901_ (.B1(net634),
    .VDD(VPWR),
    .Y(_0942_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[43] ),
    .A2(net563));
 sg13g2_a21oi_1 _2902_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1018_),
    .A2(net563),
    .Y(_0251_),
    .B1(_0942_));
 sg13g2_o21ai_1 _2903_ (.B1(net639),
    .VDD(VPWR),
    .Y(_0943_),
    .VSS(VGND),
    .A1(net693),
    .A2(net575));
 sg13g2_a21oi_1 _2904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1017_),
    .A2(net575),
    .Y(_0252_),
    .B1(_0943_));
 sg13g2_o21ai_1 _2905_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0944_),
    .VSS(VGND),
    .A1(net664),
    .A2(net574));
 sg13g2_a21oi_1 _2906_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1016_),
    .A2(net574),
    .Y(_0253_),
    .B1(_0944_));
 sg13g2_o21ai_1 _2907_ (.B1(net639),
    .VDD(VPWR),
    .Y(_0945_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[46] ),
    .A2(net574));
 sg13g2_a21oi_1 _2908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1015_),
    .A2(net574),
    .Y(_0254_),
    .B1(_0945_));
 sg13g2_o21ai_1 _2909_ (.B1(net657),
    .VDD(VPWR),
    .Y(_0946_),
    .VSS(VGND),
    .A1(net413),
    .A2(net606));
 sg13g2_a21oi_1 _2910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1014_),
    .A2(net606),
    .Y(_0255_),
    .B1(_0946_));
 sg13g2_o21ai_1 _2911_ (.B1(net657),
    .VDD(VPWR),
    .Y(_0947_),
    .VSS(VGND),
    .A1(net407),
    .A2(net609));
 sg13g2_a21oi_1 _2912_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1013_),
    .A2(net607),
    .Y(_0256_),
    .B1(_0947_));
 sg13g2_o21ai_1 _2913_ (.B1(net657),
    .VDD(VPWR),
    .Y(_0948_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[49] ),
    .A2(net610));
 sg13g2_a21oi_1 _2914_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1012_),
    .A2(net609),
    .Y(_0257_),
    .B1(_0948_));
 sg13g2_o21ai_1 _2915_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0949_),
    .VSS(VGND),
    .A1(net434),
    .A2(net608));
 sg13g2_a21oi_1 _2916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1011_),
    .A2(net608),
    .Y(_0258_),
    .B1(_0949_));
 sg13g2_o21ai_1 _2917_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0950_),
    .VSS(VGND),
    .A1(net432),
    .A2(net588));
 sg13g2_a21oi_1 _2918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1010_),
    .A2(net588),
    .Y(_0259_),
    .B1(_0950_));
 sg13g2_o21ai_1 _2919_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0951_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[52] ),
    .A2(net588));
 sg13g2_a21oi_1 _2920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1009_),
    .A2(net588),
    .Y(_0260_),
    .B1(_0951_));
 sg13g2_o21ai_1 _2921_ (.B1(net646),
    .VDD(VPWR),
    .Y(_0952_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[53] ),
    .A2(net591));
 sg13g2_a21oi_1 _2922_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1008_),
    .A2(net591),
    .Y(_0261_),
    .B1(_0952_));
 sg13g2_o21ai_1 _2923_ (.B1(net647),
    .VDD(VPWR),
    .Y(_0953_),
    .VSS(VGND),
    .A1(net726),
    .A2(net589));
 sg13g2_a21oi_1 _2924_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1007_),
    .A2(net589),
    .Y(_0262_),
    .B1(_0953_));
 sg13g2_o21ai_1 _2925_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0954_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[55] ),
    .A2(net598));
 sg13g2_a21oi_1 _2926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1006_),
    .A2(net589),
    .Y(_0263_),
    .B1(_0954_));
 sg13g2_o21ai_1 _2927_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0955_),
    .VSS(VGND),
    .A1(net804),
    .A2(net593));
 sg13g2_a21oi_1 _2928_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1005_),
    .A2(net593),
    .Y(_0264_),
    .B1(_0955_));
 sg13g2_o21ai_1 _2929_ (.B1(net644),
    .VDD(VPWR),
    .Y(_0956_),
    .VSS(VGND),
    .A1(net426),
    .A2(net587));
 sg13g2_a21oi_1 _2930_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1004_),
    .A2(net587),
    .Y(_0265_),
    .B1(_0956_));
 sg13g2_o21ai_1 _2931_ (.B1(net644),
    .VDD(VPWR),
    .Y(_0957_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[58] ),
    .A2(net583));
 sg13g2_a21oi_1 _2932_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1003_),
    .A2(net591),
    .Y(_0266_),
    .B1(_0957_));
 sg13g2_o21ai_1 _2933_ (.B1(net642),
    .VDD(VPWR),
    .Y(_0958_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[59] ),
    .A2(net582));
 sg13g2_a21oi_1 _2934_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1002_),
    .A2(net582),
    .Y(_0267_),
    .B1(_0958_));
 sg13g2_o21ai_1 _2935_ (.B1(net630),
    .VDD(VPWR),
    .Y(_0959_),
    .VSS(VGND),
    .A1(net807),
    .A2(net560));
 sg13g2_a21oi_1 _2936_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1001_),
    .A2(net560),
    .Y(_0268_),
    .B1(_0959_));
 sg13g2_o21ai_1 _2937_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0960_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[61] ),
    .A2(net556));
 sg13g2_a21oi_1 _2938_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1000_),
    .A2(net556),
    .Y(_0269_),
    .B1(_0960_));
 sg13g2_o21ai_1 _2939_ (.B1(net625),
    .VDD(VPWR),
    .Y(_0961_),
    .VSS(VGND),
    .A1(net758),
    .A2(net550));
 sg13g2_a21oi_1 _2940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0999_),
    .A2(net553),
    .Y(_0270_),
    .B1(_0961_));
 sg13g2_o21ai_1 _2941_ (.B1(net625),
    .VDD(VPWR),
    .Y(_0962_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[63] ),
    .A2(net546));
 sg13g2_a21oi_1 _2942_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0998_),
    .A2(net548),
    .Y(_0271_),
    .B1(_0962_));
 sg13g2_o21ai_1 _2943_ (.B1(net625),
    .VDD(VPWR),
    .Y(_0963_),
    .VSS(VGND),
    .A1(net328),
    .A2(net549));
 sg13g2_a21oi_1 _2944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0997_),
    .A2(net549),
    .Y(_0272_),
    .B1(_0963_));
 sg13g2_o21ai_1 _2945_ (.B1(net629),
    .VDD(VPWR),
    .Y(_0964_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[65] ),
    .A2(net552));
 sg13g2_a21oi_1 _2946_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0996_),
    .A2(net552),
    .Y(_0273_),
    .B1(_0964_));
 sg13g2_o21ai_1 _2947_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0965_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[66] ),
    .A2(net562));
 sg13g2_a21oi_1 _2948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0995_),
    .A2(net562),
    .Y(_0274_),
    .B1(_0965_));
 sg13g2_o21ai_1 _2949_ (.B1(net632),
    .VDD(VPWR),
    .Y(_0966_),
    .VSS(VGND),
    .A1(net767),
    .A2(net563));
 sg13g2_a21oi_1 _2950_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0994_),
    .A2(net563),
    .Y(_0275_),
    .B1(_0966_));
 sg13g2_o21ai_1 _2951_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0967_),
    .VSS(VGND),
    .A1(net675),
    .A2(net572));
 sg13g2_a21oi_1 _2952_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0993_),
    .A2(net572),
    .Y(_0276_),
    .B1(_0967_));
 sg13g2_o21ai_1 _2953_ (.B1(net638),
    .VDD(VPWR),
    .Y(_0968_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[69] ),
    .A2(net572));
 sg13g2_a21oi_1 _2954_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0992_),
    .A2(net572),
    .Y(_0277_),
    .B1(_0968_));
 sg13g2_o21ai_1 _2955_ (.B1(net655),
    .VDD(VPWR),
    .Y(_0969_),
    .VSS(VGND),
    .A1(net803),
    .A2(net606));
 sg13g2_a21oi_1 _2956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0991_),
    .A2(net606),
    .Y(_0278_),
    .B1(_0969_));
 sg13g2_o21ai_1 _2957_ (.B1(net656),
    .VDD(VPWR),
    .Y(_0970_),
    .VSS(VGND),
    .A1(net669),
    .A2(net609));
 sg13g2_a21oi_1 _2958_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0990_),
    .A2(net609),
    .Y(_0279_),
    .B1(_0970_));
 sg13g2_o21ai_1 _2959_ (.B1(net662),
    .VDD(VPWR),
    .Y(_0971_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[72] ),
    .A2(net617));
 sg13g2_a21oi_1 _2960_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0989_),
    .A2(net617),
    .Y(_0280_),
    .B1(_0971_));
 sg13g2_o21ai_1 _2961_ (.B1(net660),
    .VDD(VPWR),
    .Y(_0972_),
    .VSS(VGND),
    .A1(net346),
    .A2(net616));
 sg13g2_a21oi_1 _2962_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0988_),
    .A2(net616),
    .Y(_0281_),
    .B1(_0972_));
 sg13g2_o21ai_1 _2963_ (.B1(net661),
    .VDD(VPWR),
    .Y(_0973_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[74] ),
    .A2(net619));
 sg13g2_a21oi_1 _2964_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0987_),
    .A2(net619),
    .Y(_0282_),
    .B1(_0973_));
 sg13g2_o21ai_1 _2965_ (.B1(net651),
    .VDD(VPWR),
    .Y(_0974_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[75] ),
    .A2(net601));
 sg13g2_a21oi_1 _2966_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0986_),
    .A2(net620),
    .Y(_0283_),
    .B1(_0974_));
 sg13g2_o21ai_1 _2967_ (.B1(net653),
    .VDD(VPWR),
    .Y(_0975_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[76] ),
    .A2(net601));
 sg13g2_a21oi_1 _2968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0985_),
    .A2(net601),
    .Y(_0284_),
    .B1(_0975_));
 sg13g2_o21ai_1 _2969_ (.B1(net652),
    .VDD(VPWR),
    .Y(_0976_),
    .VSS(VGND),
    .A1(net826),
    .A2(net600));
 sg13g2_a21oi_1 _2970_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0984_),
    .A2(net600),
    .Y(_0285_),
    .B1(_0976_));
 sg13g2_o21ai_1 _2971_ (.B1(net649),
    .VDD(VPWR),
    .Y(_0977_),
    .VSS(VGND),
    .A1(\controller.inst_mem.mem_data[78] ),
    .A2(net595));
 sg13g2_a21oi_1 _2972_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0983_),
    .A2(net600),
    .Y(_0286_),
    .B1(_0977_));
 sg13g2_o21ai_1 _2973_ (.B1(net650),
    .VDD(VPWR),
    .Y(_0978_),
    .VSS(VGND),
    .A1(net691),
    .A2(net595));
 sg13g2_a21oi_1 _2974_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0982_),
    .A2(net595),
    .Y(_0287_),
    .B1(_0978_));
 sg13g2_o21ai_1 _2975_ (.B1(net648),
    .VDD(VPWR),
    .Y(_0979_),
    .VSS(VGND),
    .A1(net414),
    .A2(net594));
 sg13g2_a21oi_1 _2976_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0981_),
    .A2(net594),
    .Y(_0288_),
    .B1(_0979_));
 sg13g2_dfrbpq_1 _2977_ (.RESET_B(net115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net415),
    .Q(\controller.inst_mem.mem_data[81] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2978_ (.RESET_B(net168),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\controller.inst_mem.mem_data[82] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2979_ (.RESET_B(net166),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net678),
    .Q(\controller.inst_mem.mem_data[83] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2980_ (.RESET_B(net164),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\controller.inst_mem.mem_data[84] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2981_ (.RESET_B(net162),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net725),
    .Q(\controller.inst_mem.mem_data[85] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2982_ (.RESET_B(net160),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0005_),
    .Q(\controller.inst_mem.mem_data[86] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2983_ (.RESET_B(net158),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net785),
    .Q(\controller.inst_mem.mem_data[87] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2984_ (.RESET_B(net156),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0007_),
    .Q(\controller.inst_mem.mem_data[88] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2985_ (.RESET_B(net154),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net371),
    .Q(\controller.inst_mem.mem_data[89] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2986_ (.RESET_B(net152),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0009_),
    .Q(\controller.inst_mem.mem_data[90] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2987_ (.RESET_B(net150),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net424),
    .Q(\controller.inst_mem.mem_data[91] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2988_ (.RESET_B(net148),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net443),
    .Q(\controller.inst_mem.mem_data[92] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2989_ (.RESET_B(net146),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0012_),
    .Q(\controller.inst_mem.mem_data[93] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2990_ (.RESET_B(net144),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net343),
    .Q(\controller.inst_mem.mem_data[94] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2991_ (.RESET_B(net142),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net802),
    .Q(\controller.inst_mem.mem_data[95] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2992_ (.RESET_B(net140),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0015_),
    .Q(\controller.inst_mem.mem_data[96] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2993_ (.RESET_B(net138),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0016_),
    .Q(\controller.inst_mem.mem_data[97] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2994_ (.RESET_B(net136),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net422),
    .Q(\controller.inst_mem.mem_data[98] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2995_ (.RESET_B(net134),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net709),
    .Q(\controller.inst_mem.mem_data[99] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _2996_ (.RESET_B(net132),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net817),
    .Q(\controller.inst_mem.mem_data[100] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2997_ (.RESET_B(net130),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net837),
    .Q(\controller.inst_mem.mem_data[101] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _2998_ (.RESET_B(net128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net861),
    .Q(\controller.inst_mem.mem_data[102] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2999_ (.RESET_B(net126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net866),
    .Q(\controller.inst_mem.mem_data[103] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3000_ (.RESET_B(net124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0023_),
    .Q(\controller.inst_mem.mem_data[104] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3001_ (.RESET_B(net122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net389),
    .Q(\controller.inst_mem.mem_data[105] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3002_ (.RESET_B(net120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0025_),
    .Q(\controller.inst_mem.mem_data[106] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3003_ (.RESET_B(net118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net417),
    .Q(\controller.inst_mem.mem_data[107] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3004_ (.RESET_B(net116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net776),
    .Q(\controller.inst_mem.mem_data[108] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3005_ (.RESET_B(net114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0028_),
    .Q(\controller.inst_mem.mem_data[109] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3006_ (.RESET_B(net112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0029_),
    .Q(\controller.inst_mem.mem_data[110] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3007_ (.RESET_B(net110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0030_),
    .Q(\controller.inst_mem.mem_data[111] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3008_ (.RESET_B(net108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net731),
    .Q(\controller.inst_mem.mem_data[112] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3009_ (.RESET_B(net106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0032_),
    .Q(\controller.inst_mem.mem_data[113] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3010_ (.RESET_B(net104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net387),
    .Q(\controller.inst_mem.mem_data[114] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3011_ (.RESET_B(net102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net764),
    .Q(\controller.inst_mem.mem_data[115] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3012_ (.RESET_B(net100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\controller.inst_mem.mem_data[116] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3013_ (.RESET_B(net98),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net674),
    .Q(\controller.inst_mem.mem_data[117] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3014_ (.RESET_B(net96),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\controller.inst_mem.mem_data[118] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3015_ (.RESET_B(net94),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net769),
    .Q(\controller.inst_mem.mem_data[119] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3016_ (.RESET_B(net92),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\controller.inst_mem.mem_data[120] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3017_ (.RESET_B(net90),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\controller.inst_mem.mem_data[121] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3018_ (.RESET_B(net88),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\controller.inst_mem.mem_data[122] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _3019_ (.RESET_B(net86),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net363),
    .Q(\controller.inst_mem.mem_data[123] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3020_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net743),
    .Q(\controller.inst_mem.mem_data[124] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3021_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0044_),
    .Q(\controller.inst_mem.mem_data[125] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3022_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net383),
    .Q(\controller.inst_mem.mem_data[126] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3023_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net667),
    .Q(\controller.inst_mem.mem_data[127] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3024_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\controller.inst_mem.mem_data[128] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3025_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0048_),
    .Q(\controller.inst_mem.mem_data[129] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3026_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net341),
    .Q(\controller.inst_mem.mem_data[130] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3027_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net406),
    .Q(\controller.inst_mem.mem_data[131] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3028_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\controller.inst_mem.mem_data[132] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3029_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\controller.inst_mem.mem_data[133] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3030_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net385),
    .Q(\controller.inst_mem.mem_data[134] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3031_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net429),
    .Q(\controller.inst_mem.mem_data[135] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3032_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0055_),
    .Q(\controller.inst_mem.mem_data[136] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3033_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0056_),
    .Q(\controller.inst_mem.mem_data[137] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3034_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net352),
    .Q(\controller.inst_mem.mem_data[138] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3035_ (.RESET_B(net54),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net356),
    .Q(\controller.inst_mem.mem_data[139] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3036_ (.RESET_B(net52),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net412),
    .Q(\controller.inst_mem.mem_data[140] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3037_ (.RESET_B(net50),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\controller.inst_mem.mem_data[141] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3038_ (.RESET_B(net48),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net331),
    .Q(\controller.inst_mem.mem_data[142] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3039_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net369),
    .Q(\controller.inst_mem.mem_data[143] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3040_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(\controller.inst_mem.mem_data[144] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3041_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net333),
    .Q(\controller.inst_mem.mem_data[145] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3042_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net680),
    .Q(\controller.inst_mem.mem_data[146] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3043_ (.RESET_B(net327),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\controller.inst_mem.mem_data[147] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3044_ (.RESET_B(net325),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net437),
    .Q(\controller.inst_mem.mem_data[148] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3045_ (.RESET_B(net323),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\controller.inst_mem.mem_data[149] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3046_ (.RESET_B(net321),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\controller.inst_mem.mem_data[150] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3047_ (.RESET_B(net319),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net358),
    .Q(\controller.inst_mem.mem_data[151] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3048_ (.RESET_B(net317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\controller.inst_mem.mem_data[152] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3049_ (.RESET_B(net315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net772),
    .Q(\controller.inst_mem.mem_data[153] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3050_ (.RESET_B(net313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\controller.inst_mem.mem_data[154] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3051_ (.RESET_B(net311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\controller.inst_mem.mem_data[155] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3052_ (.RESET_B(net309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net704),
    .Q(\controller.inst_mem.mem_data[156] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3053_ (.RESET_B(net307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\controller.inst_mem.mem_data[157] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3054_ (.RESET_B(net305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\controller.inst_mem.mem_data[158] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3055_ (.RESET_B(net303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net795),
    .Q(\controller.inst_mem.mem_data[159] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3056_ (.RESET_B(net301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\controller.inst_mem.mem_data[160] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3057_ (.RESET_B(net299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\controller.inst_mem.mem_data[161] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3058_ (.RESET_B(net297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net339),
    .Q(\controller.inst_mem.mem_data[162] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3059_ (.RESET_B(net295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\controller.inst_mem.mem_data[163] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3060_ (.RESET_B(net293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\controller.inst_mem.mem_data[164] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3061_ (.RESET_B(net291),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\controller.inst_mem.mem_data[165] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3062_ (.RESET_B(net289),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net360),
    .Q(\controller.inst_mem.mem_data[166] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3063_ (.RESET_B(net287),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\controller.inst_mem.mem_data[167] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3064_ (.RESET_B(net285),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\controller.inst_mem.mem_data[168] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3065_ (.RESET_B(net283),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net337),
    .Q(\controller.inst_mem.mem_data[169] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3066_ (.RESET_B(net281),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net754),
    .Q(\controller.inst_mem.mem_data[170] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3067_ (.RESET_B(net279),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0090_),
    .Q(\controller.inst_mem.mem_data[171] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3068_ (.RESET_B(net277),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net745),
    .Q(\controller.inst_mem.mem_data[172] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3069_ (.RESET_B(net275),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\controller.inst_mem.mem_data[173] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3070_ (.RESET_B(net273),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\controller.inst_mem.mem_data[174] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3071_ (.RESET_B(net271),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\controller.inst_mem.mem_data[175] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3072_ (.RESET_B(net269),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net700),
    .Q(\controller.inst_mem.mem_data[176] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3073_ (.RESET_B(net267),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\controller.inst_mem.mem_data[177] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3074_ (.RESET_B(net265),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net698),
    .Q(\controller.inst_mem.mem_data[178] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _3075_ (.RESET_B(net263),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\controller.inst_mem.mem_data[179] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3076_ (.RESET_B(net261),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\controller.inst_mem.mem_data[180] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3077_ (.RESET_B(net259),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net399),
    .Q(\controller.inst_mem.mem_data[181] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3078_ (.RESET_B(net257),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net849),
    .Q(\controller.inst_mem.mem_data[182] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3079_ (.RESET_B(net255),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\controller.inst_mem.mem_data[183] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3080_ (.RESET_B(net253),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net379),
    .Q(\controller.inst_mem.mem_data[184] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3081_ (.RESET_B(net251),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\controller.inst_mem.mem_data[185] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3082_ (.RESET_B(net249),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net431),
    .Q(\controller.inst_mem.mem_data[186] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3083_ (.RESET_B(net247),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net815),
    .Q(\controller.inst_mem.mem_data[187] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3084_ (.RESET_B(net245),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\controller.inst_mem.mem_data[188] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3085_ (.RESET_B(net243),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net439),
    .Q(\controller.inst_mem.mem_data[189] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3086_ (.RESET_B(net241),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\controller.inst_mem.mem_data[190] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3087_ (.RESET_B(net239),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net381),
    .Q(\controller.inst_mem.mem_data[191] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3088_ (.RESET_B(net237),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net395),
    .Q(\controller.inst_mem.mem_data[192] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3089_ (.RESET_B(net235),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\controller.inst_mem.mem_data[193] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3090_ (.RESET_B(net233),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0113_),
    .Q(\controller.inst_mem.mem_data[194] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _3091_ (.RESET_B(net231),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net401),
    .Q(\controller.inst_mem.mem_data[195] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3092_ (.RESET_B(net229),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net791),
    .Q(\controller.inst_mem.mem_data[196] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3093_ (.RESET_B(net227),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\controller.inst_mem.mem_data[197] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3094_ (.RESET_B(net225),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net712),
    .Q(\controller.inst_mem.mem_data[198] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _3095_ (.RESET_B(net223),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net756),
    .Q(\controller.inst_mem.mem_data[199] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3096_ (.RESET_B(net221),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net830),
    .Q(\controller.extended_jump_target[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3097_ (.RESET_B(net219),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net845),
    .Q(\controller.extended_jump_target[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _3098_ (.RESET_B(net217),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\controller.extended_jump_target[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3099_ (.RESET_B(net215),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\controller.inst_mem.extended_word[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3100_ (.RESET_B(net213),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\controller.inst_mem.extended_word[4] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3101_ (.RESET_B(net211),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net335),
    .Q(\controller.inst_mem.extended_word[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3102_ (.RESET_B(net209),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\controller.inst_mem.extended_word[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3103_ (.RESET_B(net207),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net702),
    .Q(\controller.inst_mem.extended_word[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3104_ (.RESET_B(net205),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\controller.inst_mem.extended_word[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _3105_ (.RESET_B(net203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net762),
    .Q(\controller.extended_cond.opcode[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _3106_ (.RESET_B(net201),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net937),
    .Q(\controller.extended_cond.opcode[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3107_ (.RESET_B(net199),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\controller.extended_cond.opcode[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3108_ (.RESET_B(net197),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\controller.extended_then_action[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3109_ (.RESET_B(net195),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\controller.extended_then_action[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _3110_ (.RESET_B(net193),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\controller.extended_then_action[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3111_ (.RESET_B(net191),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net686),
    .Q(\controller.extended_then_action[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3112_ (.RESET_B(net189),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\controller.extended_then_action[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3113_ (.RESET_B(net187),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\controller.extended_then_action[5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3114_ (.RESET_B(net185),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\controller.inst_mem.extended_word[18] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3115_ (.RESET_B(net183),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net365),
    .Q(\controller.inst_mem.extended_word[19] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3116_ (.RESET_B(net181),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net393),
    .Q(\controller.inst_mem.extended_word[20] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3117_ (.RESET_B(net179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net404),
    .Q(\controller.inst_mem.extended_word[21] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3118_ (.RESET_B(net177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\controller.inst_mem.extended_word[22] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3119_ (.RESET_B(net175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net354),
    .Q(\controller.inst_mem.extended_word[23] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3120_ (.RESET_B(net173),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\controller.extended_state[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3121_ (.RESET_B(net171),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net377),
    .Q(\controller.extended_state[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3122_ (.RESET_B(net169),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net752),
    .Q(\controller.extended_state[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3123_ (.RESET_B(net165),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\controller.inst_mem.addr[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _3124_ (.RESET_B(net161),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net979),
    .Q(\controller.inst_mem.addr[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3125_ (.RESET_B(net157),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net987),
    .Q(\controller.inst_mem.addr[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _3126_ (.RESET_B(net153),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net968),
    .Q(\controller.alu_buffer.buffer[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3127_ (.RESET_B(net149),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net972),
    .Q(\controller.alu_buffer.buffer[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3128_ (.RESET_B(net145),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\controller.alu_buffer.buffer[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3129_ (.RESET_B(net141),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\controller.alu_buffer.buffer[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3130_ (.RESET_B(net137),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\controller.alu_buffer.buffer[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3131_ (.RESET_B(net133),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net981),
    .Q(\controller.alu_buffer.buffer[4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3132_ (.RESET_B(net129),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net962),
    .Q(\controller.alu_buffer.buffer[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3133_ (.RESET_B(net125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\controller.alu_buffer.buffer[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _3134_ (.RESET_B(net121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net974),
    .Q(\controller.alu_buffer.buffer[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3135_ (.RESET_B(net117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net964),
    .Q(\controller.alu_buffer.buffer[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3136_ (.RESET_B(net113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net935),
    .Q(\controller.alu_buffer.buffer[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3137_ (.RESET_B(net109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net976),
    .Q(\controller.alu_buffer.buffer[11] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3138_ (.RESET_B(net105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net970),
    .Q(\controller.alu_buffer.buffer[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3139_ (.RESET_B(net101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net955),
    .Q(\controller.alu_buffer.buffer[13] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3140_ (.RESET_B(net97),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net951),
    .Q(\controller.alu_buffer.buffer[14] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3141_ (.RESET_B(net93),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net923),
    .Q(\controller.alu_buffer.buffer[15] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3142_ (.RESET_B(net89),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net966),
    .Q(\controller.alu_buffer.buffer[16] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _3143_ (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net959),
    .Q(\controller.alu_buffer.buffer[17] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _3144_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net953),
    .Q(\controller.alu_buffer.buffer[18] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _3145_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net946),
    .Q(\controller.alu_buffer.buffer[19] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _3146_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net949),
    .Q(\controller.alu_buffer.buffer[20] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _3147_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\controller.alu_buffer.buffer[21] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _3148_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net957),
    .Q(\controller.alu_buffer.buffer[22] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3149_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net914),
    .Q(\controller.alu_buffer.buffer[23] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3150_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\controller.output_controller.keep[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3151_ (.RESET_B(net55),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net941),
    .Q(\controller.output_controller.keep[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3152_ (.RESET_B(net53),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net918),
    .Q(\controller.output_controller.keep[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _3153_ (.RESET_B(net51),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\controller.counter2.counter_0[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3154_ (.RESET_B(net47),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net931),
    .Q(\controller.counter2.counter_0[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3155_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net920),
    .Q(\controller.counter2.counter_0[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3156_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net929),
    .Q(\controller.counter2.counter_0[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3157_ (.RESET_B(net324),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\controller.counter2.counter_0[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _3158_ (.RESET_B(net320),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net939),
    .Q(\controller.counter2.counter_0[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3159_ (.RESET_B(net316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net895),
    .Q(\controller.counter2.counter_0[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3160_ (.RESET_B(net312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net880),
    .Q(\controller.counter2.counter_0[7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _3161_ (.RESET_B(net308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\controller.counter2.counter_0[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3162_ (.RESET_B(net304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net887),
    .Q(\controller.counter2.counter_0[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3163_ (.RESET_B(net300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net925),
    .Q(\controller.counter2.counter_0[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _3164_ (.RESET_B(net296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net898),
    .Q(\controller.counter2.counter_0[11] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _3165_ (.RESET_B(net292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0188_),
    .Q(\controller.counter2.counter_0[12] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3166_ (.RESET_B(net288),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net900),
    .Q(\controller.counter2.counter_0[13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _3167_ (.RESET_B(net284),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\controller.counter2.counter_0[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3168_ (.RESET_B(net280),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\controller.counter2.counter_0[15] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3169_ (.RESET_B(net276),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\controller.counter2.counter_1[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _3170_ (.RESET_B(net272),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\controller.counter2.counter_1[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3171_ (.RESET_B(net268),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net912),
    .Q(\controller.counter2.counter_1[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3172_ (.RESET_B(net264),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net891),
    .Q(\controller.counter2.counter_1[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _3173_ (.RESET_B(net260),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0196_),
    .Q(\controller.counter2.counter_1[4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3174_ (.RESET_B(net256),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0197_),
    .Q(\controller.counter2.counter_1[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3175_ (.RESET_B(net252),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net889),
    .Q(\controller.counter2.counter_1[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _3176_ (.RESET_B(net248),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0199_),
    .Q(\controller.counter2.counter_1[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3177_ (.RESET_B(net244),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0200_),
    .Q(\controller.counter2.counter_1[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3178_ (.RESET_B(net240),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net902),
    .Q(\controller.counter2.counter_1[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3179_ (.RESET_B(net236),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net908),
    .Q(\controller.counter2.counter_1[10] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3180_ (.RESET_B(net232),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net884),
    .Q(\controller.counter2.counter_1[11] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _3181_ (.RESET_B(net228),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0204_),
    .Q(\controller.counter2.counter_1[12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _3182_ (.RESET_B(net224),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net927),
    .Q(\controller.counter2.counter_1[13] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3183_ (.RESET_B(net220),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net905),
    .Q(\controller.counter2.counter_1[14] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3184_ (.RESET_B(net216),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\controller.counter2.counter_1[15] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3185_ (.RESET_B(net212),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0208_),
    .Q(\controller.const_data[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3186_ (.RESET_B(net208),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net672),
    .Q(\controller.const_data[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3187_ (.RESET_B(net204),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net696),
    .Q(\controller.const_data[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3188_ (.RESET_B(net200),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net833),
    .Q(\controller.const_data[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3189_ (.RESET_B(net196),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0212_),
    .Q(\controller.const_data[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3190_ (.RESET_B(net192),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net420),
    .Q(\controller.const_data[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3191_ (.RESET_B(net188),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0214_),
    .Q(\controller.const_data[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3192_ (.RESET_B(net184),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net716),
    .Q(\controller.const_data[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3193_ (.RESET_B(net180),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0216_),
    .Q(\controller.const_data[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3194_ (.RESET_B(net176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0217_),
    .Q(\controller.const_data[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3195_ (.RESET_B(net172),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net391),
    .Q(\controller.const_data[10] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3196_ (.RESET_B(net167),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0219_),
    .Q(\controller.const_data[11] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3197_ (.RESET_B(net159),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0220_),
    .Q(\controller.const_data[12] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3198_ (.RESET_B(net151),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net373),
    .Q(\controller.const_data[13] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3199_ (.RESET_B(net143),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\controller.const_data[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _3200_ (.RESET_B(net135),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\controller.const_data[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3201_ (.RESET_B(net127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net349),
    .Q(\controller.const_data[16] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3202_ (.RESET_B(net119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0225_),
    .Q(\controller.const_data[17] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3203_ (.RESET_B(net111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\controller.const_data[18] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3204_ (.RESET_B(net103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\controller.const_data[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3205_ (.RESET_B(net95),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net345),
    .Q(\controller.const_data[20] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3206_ (.RESET_B(net87),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0229_),
    .Q(\controller.const_data[21] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3207_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net719),
    .Q(\controller.const_data[22] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3208_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0231_),
    .Q(\controller.const_data[23] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3209_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0232_),
    .Q(\controller.const_data[24] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3210_ (.RESET_B(net49),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0233_),
    .Q(\controller.const_data[25] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _3211_ (.RESET_B(net41),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net688),
    .Q(\controller.const_data[26] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3212_ (.RESET_B(net322),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0235_),
    .Q(\controller.const_data[27] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3213_ (.RESET_B(net314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net397),
    .Q(\controller.const_data[28] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3214_ (.RESET_B(net306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0237_),
    .Q(\controller.const_data[29] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3215_ (.RESET_B(net298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net441),
    .Q(\controller.const_data[30] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3216_ (.RESET_B(net290),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net690),
    .Q(\controller.const_data[31] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3217_ (.RESET_B(net282),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0240_),
    .Q(\controller.inst_mem.mem_data[32] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3218_ (.RESET_B(net274),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\controller.inst_mem.mem_data[33] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3219_ (.RESET_B(net266),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net721),
    .Q(\controller.inst_mem.mem_data[34] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3220_ (.RESET_B(net258),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0243_),
    .Q(\controller.inst_mem.mem_data[35] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3221_ (.RESET_B(net250),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net749),
    .Q(\controller.inst_mem.mem_data[36] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3222_ (.RESET_B(net242),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\controller.inst_mem.mem_data[37] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3223_ (.RESET_B(net234),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net870),
    .Q(\controller.inst_mem.mem_data[38] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3224_ (.RESET_B(net226),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0247_),
    .Q(\controller.inst_mem.mem_data[39] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3225_ (.RESET_B(net218),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0248_),
    .Q(\controller.inst_mem.mem_data[40] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3226_ (.RESET_B(net210),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net723),
    .Q(\controller.inst_mem.mem_data[41] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3227_ (.RESET_B(net202),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0250_),
    .Q(\controller.inst_mem.mem_data[42] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3228_ (.RESET_B(net194),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net741),
    .Q(\controller.inst_mem.mem_data[43] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3229_ (.RESET_B(net186),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0252_),
    .Q(\controller.inst_mem.mem_data[44] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3230_ (.RESET_B(net178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0253_),
    .Q(\controller.inst_mem.mem_data[45] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3231_ (.RESET_B(net170),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net665),
    .Q(\controller.inst_mem.mem_data[46] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3232_ (.RESET_B(net155),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0255_),
    .Q(\controller.inst_mem.mem_data[47] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3233_ (.RESET_B(net139),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\controller.inst_mem.mem_data[48] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3234_ (.RESET_B(net123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net408),
    .Q(\controller.inst_mem.mem_data[49] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3235_ (.RESET_B(net107),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0258_),
    .Q(\controller.inst_mem.mem_data[50] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3236_ (.RESET_B(net91),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0259_),
    .Q(\controller.inst_mem.mem_data[51] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3237_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net433),
    .Q(\controller.inst_mem.mem_data[52] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3238_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net787),
    .Q(\controller.inst_mem.mem_data[53] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3239_ (.RESET_B(net326),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0262_),
    .Q(\controller.inst_mem.mem_data[54] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3240_ (.RESET_B(net310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net727),
    .Q(\controller.inst_mem.mem_data[55] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3241_ (.RESET_B(net294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\controller.inst_mem.mem_data[56] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3242_ (.RESET_B(net278),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0265_),
    .Q(\controller.inst_mem.mem_data[57] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3243_ (.RESET_B(net262),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net427),
    .Q(\controller.inst_mem.mem_data[58] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3244_ (.RESET_B(net246),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net766),
    .Q(\controller.inst_mem.mem_data[59] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3245_ (.RESET_B(net230),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0268_),
    .Q(\controller.inst_mem.mem_data[60] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3246_ (.RESET_B(net214),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net808),
    .Q(\controller.inst_mem.mem_data[61] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3247_ (.RESET_B(net198),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0270_),
    .Q(\controller.inst_mem.mem_data[62] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3248_ (.RESET_B(net182),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net759),
    .Q(\controller.inst_mem.mem_data[63] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3249_ (.RESET_B(net163),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0272_),
    .Q(\controller.inst_mem.mem_data[64] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3250_ (.RESET_B(net131),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net329),
    .Q(\controller.inst_mem.mem_data[65] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3251_ (.RESET_B(net99),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net375),
    .Q(\controller.inst_mem.mem_data[66] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3252_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0275_),
    .Q(\controller.inst_mem.mem_data[67] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3253_ (.RESET_B(net318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0276_),
    .Q(\controller.inst_mem.mem_data[68] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3254_ (.RESET_B(net286),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net676),
    .Q(\controller.inst_mem.mem_data[69] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3255_ (.RESET_B(net254),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0278_),
    .Q(\controller.inst_mem.mem_data[70] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3256_ (.RESET_B(net222),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0279_),
    .Q(\controller.inst_mem.mem_data[71] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3257_ (.RESET_B(net190),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net670),
    .Q(\controller.inst_mem.mem_data[72] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3258_ (.RESET_B(net147),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0281_),
    .Q(\controller.inst_mem.mem_data[73] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3259_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net347),
    .Q(\controller.inst_mem.mem_data[74] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _3260_ (.RESET_B(net302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net367),
    .Q(\controller.inst_mem.mem_data[75] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3261_ (.RESET_B(net238),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net793),
    .Q(\controller.inst_mem.mem_data[76] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _3262_ (.RESET_B(net174),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0285_),
    .Q(\controller.inst_mem.mem_data[77] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3263_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net827),
    .Q(\controller.inst_mem.mem_data[78] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3264_ (.RESET_B(net206),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0287_),
    .Q(\controller.inst_mem.mem_data[79] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3265_ (.RESET_B(net270),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0288_),
    .Q(\controller.inst_mem.mem_data[80] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_tiehi _3042__40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi _3211__41 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi _3041__42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi _3155__43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi _3040__44 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi _3263__45 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi _3039__46 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi _3154__47 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi _3038__48 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi _3210__49 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi _3037__50 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi _3153__51 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi _3036__52 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi _3152__53 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi _3035__54 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi _3151__55 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_tiehi _3034__56 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi _3150__57 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi _3033__58 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi _3238__59 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi _3032__60 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi _3149__61 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi _3031__62 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi _3209__63 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi _3030__64 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi _3148__65 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi _3029__66 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi _3252__67 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi _3028__68 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi _3147__69 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi _3027__70 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi _3208__71 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi _3026__72 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi _3146__73 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi _3025__74 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi _3237__75 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_tiehi _3024__76 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net76));
 sg13g2_tiehi _3145__77 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net77));
 sg13g2_tiehi _3023__78 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net78));
 sg13g2_tiehi _3207__79 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net79));
 sg13g2_tiehi _3022__80 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net80));
 sg13g2_tiehi _3144__81 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net81));
 sg13g2_tiehi _3021__82 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net82));
 sg13g2_tiehi _3259__83 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net83));
 sg13g2_tiehi _3020__84 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net84));
 sg13g2_tiehi _3143__85 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net85));
 sg13g2_tiehi _3019__86 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net86));
 sg13g2_tiehi _3206__87 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net87));
 sg13g2_tiehi _3018__88 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net88));
 sg13g2_tiehi _3142__89 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net89));
 sg13g2_tiehi _3017__90 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net90));
 sg13g2_tiehi _3236__91 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net91));
 sg13g2_tiehi _3016__92 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net92));
 sg13g2_tiehi _3141__93 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net93));
 sg13g2_tiehi _3015__94 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net94));
 sg13g2_tiehi _3205__95 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net95));
 sg13g2_tiehi _3014__96 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net96));
 sg13g2_tiehi _3140__97 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net97));
 sg13g2_tiehi _3013__98 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net98));
 sg13g2_tiehi _3251__99 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net99));
 sg13g2_tiehi _3012__100 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net100));
 sg13g2_tiehi _3139__101 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net101));
 sg13g2_tiehi _3011__102 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net102));
 sg13g2_tiehi _3204__103 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net103));
 sg13g2_tiehi _3010__104 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net104));
 sg13g2_tiehi _3138__105 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net105));
 sg13g2_tiehi _3009__106 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net106));
 sg13g2_tiehi _3235__107 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net107));
 sg13g2_tiehi _3008__108 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net108));
 sg13g2_tiehi _3137__109 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net109));
 sg13g2_tiehi _3007__110 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net110));
 sg13g2_tiehi _3203__111 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net111));
 sg13g2_tiehi _3006__112 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net112));
 sg13g2_tiehi _3136__113 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net113));
 sg13g2_tiehi _3005__114 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net114));
 sg13g2_tiehi _2977__115 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net115));
 sg13g2_tiehi _3004__116 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net116));
 sg13g2_tiehi _3135__117 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net117));
 sg13g2_tiehi _3003__118 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net118));
 sg13g2_tiehi _3202__119 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net119));
 sg13g2_tiehi _3002__120 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net120));
 sg13g2_tiehi _3134__121 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net121));
 sg13g2_tiehi _3001__122 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net122));
 sg13g2_tiehi _3234__123 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net123));
 sg13g2_tiehi _3000__124 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net124));
 sg13g2_tiehi _3133__125 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net125));
 sg13g2_tiehi _2999__126 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net126));
 sg13g2_tiehi _3201__127 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net127));
 sg13g2_tiehi _2998__128 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net128));
 sg13g2_tiehi _3132__129 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net129));
 sg13g2_tiehi _2997__130 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net130));
 sg13g2_tiehi _3250__131 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net131));
 sg13g2_tiehi _2996__132 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net132));
 sg13g2_tiehi _3131__133 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net133));
 sg13g2_tiehi _2995__134 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net134));
 sg13g2_tiehi _3200__135 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net135));
 sg13g2_tiehi _2994__136 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net136));
 sg13g2_tiehi _3130__137 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net137));
 sg13g2_tiehi _2993__138 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net138));
 sg13g2_tiehi _3233__139 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net139));
 sg13g2_tiehi _2992__140 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net140));
 sg13g2_tiehi _3129__141 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net141));
 sg13g2_tiehi _2991__142 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net142));
 sg13g2_tiehi _3199__143 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net143));
 sg13g2_tiehi _2990__144 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net144));
 sg13g2_tiehi _3128__145 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net145));
 sg13g2_tiehi _2989__146 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net146));
 sg13g2_tiehi _3258__147 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net147));
 sg13g2_tiehi _2988__148 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net148));
 sg13g2_tiehi _3127__149 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net149));
 sg13g2_tiehi _2987__150 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net150));
 sg13g2_tiehi _3198__151 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net151));
 sg13g2_tiehi _2986__152 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net152));
 sg13g2_tiehi _3126__153 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net153));
 sg13g2_tiehi _2985__154 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net154));
 sg13g2_tiehi _3232__155 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net155));
 sg13g2_tiehi _2984__156 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net156));
 sg13g2_tiehi _3125__157 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net157));
 sg13g2_tiehi _2983__158 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net158));
 sg13g2_tiehi _3197__159 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net159));
 sg13g2_tiehi _2982__160 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net160));
 sg13g2_tiehi _3124__161 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net161));
 sg13g2_tiehi _2981__162 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net162));
 sg13g2_tiehi _3249__163 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net163));
 sg13g2_tiehi _2980__164 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net164));
 sg13g2_tiehi _3123__165 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net165));
 sg13g2_tiehi _2979__166 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net166));
 sg13g2_tiehi _3196__167 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net167));
 sg13g2_tiehi _2978__168 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net168));
 sg13g2_tiehi _3122__169 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net169));
 sg13g2_tiehi _3231__170 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net170));
 sg13g2_tiehi _3121__171 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net171));
 sg13g2_tiehi _3195__172 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net172));
 sg13g2_tiehi _3120__173 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net173));
 sg13g2_tiehi _3262__174 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net174));
 sg13g2_tiehi _3119__175 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net175));
 sg13g2_tiehi _3194__176 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net176));
 sg13g2_tiehi _3118__177 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net177));
 sg13g2_tiehi _3230__178 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net178));
 sg13g2_tiehi _3117__179 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net179));
 sg13g2_tiehi _3193__180 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net180));
 sg13g2_tiehi _3116__181 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net181));
 sg13g2_tiehi _3248__182 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net182));
 sg13g2_tiehi _3115__183 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net183));
 sg13g2_tiehi _3192__184 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net184));
 sg13g2_tiehi _3114__185 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net185));
 sg13g2_tiehi _3229__186 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net186));
 sg13g2_tiehi _3113__187 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net187));
 sg13g2_tiehi _3191__188 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net188));
 sg13g2_tiehi _3112__189 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net189));
 sg13g2_tiehi _3257__190 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net190));
 sg13g2_tiehi _3111__191 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net191));
 sg13g2_tiehi _3190__192 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net192));
 sg13g2_tiehi _3110__193 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net193));
 sg13g2_tiehi _3228__194 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net194));
 sg13g2_tiehi _3109__195 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net195));
 sg13g2_tiehi _3189__196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net196));
 sg13g2_tiehi _3108__197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net197));
 sg13g2_tiehi _3247__198 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net198));
 sg13g2_tiehi _3107__199 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net199));
 sg13g2_tiehi _3188__200 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net200));
 sg13g2_tiehi _3106__201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net201));
 sg13g2_tiehi _3227__202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net202));
 sg13g2_tiehi _3105__203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net203));
 sg13g2_tiehi _3187__204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net204));
 sg13g2_tiehi _3104__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net205));
 sg13g2_tiehi _3264__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net206));
 sg13g2_tiehi _3103__207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net207));
 sg13g2_tiehi _3186__208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net208));
 sg13g2_tiehi _3102__209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net209));
 sg13g2_tiehi _3226__210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net210));
 sg13g2_tiehi _3101__211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net211));
 sg13g2_tiehi _3185__212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net212));
 sg13g2_tiehi _3100__213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net213));
 sg13g2_tiehi _3246__214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net214));
 sg13g2_tiehi _3099__215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net215));
 sg13g2_tiehi _3184__216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net216));
 sg13g2_tiehi _3098__217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net217));
 sg13g2_tiehi _3225__218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net218));
 sg13g2_tiehi _3097__219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_tiehi _3183__220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_tiehi _3096__221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net221));
 sg13g2_tiehi _3256__222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net222));
 sg13g2_tiehi _3095__223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net223));
 sg13g2_tiehi _3182__224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net224));
 sg13g2_tiehi _3094__225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net225));
 sg13g2_tiehi _3224__226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net226));
 sg13g2_tiehi _3093__227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net227));
 sg13g2_tiehi _3181__228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_tiehi _3092__229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_tiehi _3245__230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net230));
 sg13g2_tiehi _3091__231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net231));
 sg13g2_tiehi _3180__232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net232));
 sg13g2_tiehi _3090__233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net233));
 sg13g2_tiehi _3223__234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net234));
 sg13g2_tiehi _3089__235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net235));
 sg13g2_tiehi _3179__236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net236));
 sg13g2_tiehi _3088__237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net237));
 sg13g2_tiehi _3261__238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net238));
 sg13g2_tiehi _3087__239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net239));
 sg13g2_tiehi _3178__240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net240));
 sg13g2_tiehi _3086__241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net241));
 sg13g2_tiehi _3222__242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net242));
 sg13g2_tiehi _3085__243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net243));
 sg13g2_tiehi _3177__244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net244));
 sg13g2_tiehi _3084__245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net245));
 sg13g2_tiehi _3244__246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net246));
 sg13g2_tiehi _3083__247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net247));
 sg13g2_tiehi _3176__248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net248));
 sg13g2_tiehi _3082__249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net249));
 sg13g2_tiehi _3221__250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net250));
 sg13g2_tiehi _3081__251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net251));
 sg13g2_tiehi _3175__252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net252));
 sg13g2_tiehi _3080__253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net253));
 sg13g2_tiehi _3255__254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net254));
 sg13g2_tiehi _3079__255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net255));
 sg13g2_tiehi _3174__256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net256));
 sg13g2_tiehi _3078__257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net257));
 sg13g2_tiehi _3220__258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net258));
 sg13g2_tiehi _3077__259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net259));
 sg13g2_tiehi _3173__260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net260));
 sg13g2_tiehi _3076__261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net261));
 sg13g2_tiehi _3243__262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net262));
 sg13g2_tiehi _3075__263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net263));
 sg13g2_tiehi _3172__264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net264));
 sg13g2_tiehi _3074__265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net265));
 sg13g2_tiehi _3219__266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net266));
 sg13g2_tiehi _3073__267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net267));
 sg13g2_tiehi _3171__268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net268));
 sg13g2_tiehi _3072__269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net269));
 sg13g2_tiehi _3265__270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net270));
 sg13g2_tiehi _3071__271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net271));
 sg13g2_tiehi _3170__272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net272));
 sg13g2_tiehi _3070__273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net273));
 sg13g2_tiehi _3218__274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net274));
 sg13g2_tiehi _3069__275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net275));
 sg13g2_tiehi _3169__276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net276));
 sg13g2_tiehi _3068__277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net277));
 sg13g2_tiehi _3242__278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net278));
 sg13g2_tiehi _3067__279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net279));
 sg13g2_tiehi _3168__280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net280));
 sg13g2_tiehi _3066__281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net281));
 sg13g2_tiehi _3217__282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net282));
 sg13g2_tiehi _3065__283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net283));
 sg13g2_tiehi _3167__284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net284));
 sg13g2_tiehi _3064__285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net285));
 sg13g2_tiehi _3254__286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net286));
 sg13g2_tiehi _3063__287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net287));
 sg13g2_tiehi _3166__288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net288));
 sg13g2_tiehi _3062__289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net289));
 sg13g2_tiehi _3216__290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net290));
 sg13g2_tiehi _3061__291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net291));
 sg13g2_tiehi _3165__292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net292));
 sg13g2_tiehi _3060__293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net293));
 sg13g2_tiehi _3241__294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net294));
 sg13g2_tiehi _3059__295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net295));
 sg13g2_tiehi _3164__296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net296));
 sg13g2_tiehi _3058__297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net297));
 sg13g2_tiehi _3215__298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net298));
 sg13g2_tiehi _3057__299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net299));
 sg13g2_tiehi _3163__300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net300));
 sg13g2_tiehi _3056__301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net301));
 sg13g2_tiehi _3260__302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net302));
 sg13g2_tiehi _3055__303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net303));
 sg13g2_tiehi _3162__304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net304));
 sg13g2_tiehi _3054__305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net305));
 sg13g2_tiehi _3214__306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net306));
 sg13g2_tiehi _3053__307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net307));
 sg13g2_tiehi _3161__308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net308));
 sg13g2_tiehi _3052__309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net309));
 sg13g2_tiehi _3240__310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net310));
 sg13g2_tiehi _3051__311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net311));
 sg13g2_tiehi _3160__312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net312));
 sg13g2_tiehi _3050__313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net313));
 sg13g2_tiehi _3213__314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net314));
 sg13g2_tiehi _3049__315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net315));
 sg13g2_tiehi _3159__316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net316));
 sg13g2_tiehi _3048__317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net317));
 sg13g2_tiehi _3253__318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net318));
 sg13g2_tiehi _3047__319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net319));
 sg13g2_tiehi _3158__320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net320));
 sg13g2_tiehi _3046__321 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net321));
 sg13g2_tiehi _3212__322 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net322));
 sg13g2_tiehi _3045__323 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net323));
 sg13g2_tiehi _3157__324 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net324));
 sg13g2_tiehi _3044__325 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net325));
 sg13g2_tiehi _3239__326 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net326));
 sg13g2_tiehi _3043__327 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net327));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_can_lehmann_fsm_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net24));
 sg13g2_tielo heichips25_can_lehmann_fsm_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_tielo heichips25_can_lehmann_fsm_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo heichips25_can_lehmann_fsm_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo heichips25_can_lehmann_fsm_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo heichips25_can_lehmann_fsm_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tielo heichips25_can_lehmann_fsm_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net30));
 sg13g2_tielo heichips25_can_lehmann_fsm_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net31));
 sg13g2_tielo heichips25_can_lehmann_fsm_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_tielo heichips25_can_lehmann_fsm_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_tielo heichips25_can_lehmann_fsm_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_tielo heichips25_can_lehmann_fsm_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_tielo heichips25_can_lehmann_fsm_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_tielo heichips25_can_lehmann_fsm_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net37));
 sg13g2_tielo heichips25_can_lehmann_fsm_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net38));
 sg13g2_tiehi _3156__39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_buf_8 fanout444 (.A(net445),
    .X(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout445 (.A(_0773_),
    .X(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout446 (.A(net447),
    .X(net446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout447 (.A(_0772_),
    .X(net447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout448 (.A(net449),
    .X(net448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout449 (.A(_0770_),
    .X(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout450 (.A(net451),
    .X(net450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout451 (.A(net454),
    .X(net451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout452 (.A(net453),
    .X(net452),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout453 (.A(net454),
    .X(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout454 (.A(_0830_),
    .X(net454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout455 (.A(net456),
    .X(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout456 (.A(net457),
    .X(net456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout457 (.A(_0607_),
    .X(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout458 (.A(net459),
    .X(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout459 (.A(_0596_),
    .X(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout460 (.A(_0596_),
    .X(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout461 (.A(net465),
    .X(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout462 (.A(net465),
    .X(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout463 (.A(net465),
    .X(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout464 (.A(net465),
    .X(net464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout465 (.A(_0595_),
    .X(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout466 (.A(net467),
    .X(net466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout467 (.A(net469),
    .X(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout468 (.A(net469),
    .X(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout469 (.A(_0586_),
    .X(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout470 (.A(net473),
    .X(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout471 (.A(net473),
    .X(net471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout472 (.A(net473),
    .X(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout473 (.A(_0584_),
    .X(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout474 (.A(net475),
    .X(net474),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout475 (.A(_0748_),
    .X(net475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout476 (.A(net477),
    .X(net476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout477 (.A(net478),
    .X(net477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout478 (.A(_0748_),
    .X(net478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout479 (.A(net480),
    .X(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout480 (.A(_0731_),
    .X(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout481 (.A(net484),
    .X(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout482 (.A(net484),
    .X(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout483 (.A(net484),
    .X(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout484 (.A(_0603_),
    .X(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout485 (.A(_0545_),
    .X(net485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout486 (.A(_0474_),
    .X(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout487 (.A(_0474_),
    .X(net487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout488 (.A(_0439_),
    .X(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout489 (.A(_0438_),
    .X(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout490 (.A(_0422_),
    .X(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout491 (.A(net493),
    .X(net491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout492 (.A(net493),
    .X(net492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout493 (.A(_1232_),
    .X(net493),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout494 (.A(net497),
    .X(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout495 (.A(net497),
    .X(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout497 (.A(_1227_),
    .X(net497),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout498 (.A(net501),
    .X(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout499 (.A(net501),
    .X(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout500 (.A(net501),
    .X(net500),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout501 (.A(_1226_),
    .X(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout502 (.A(net505),
    .X(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout503 (.A(net505),
    .X(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout504 (.A(net505),
    .X(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout505 (.A(_1222_),
    .X(net505),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout506 (.A(net509),
    .X(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout507 (.A(net509),
    .X(net507),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout509 (.A(_1220_),
    .X(net509),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout510 (.A(net513),
    .X(net510),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout511 (.A(net513),
    .X(net511),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout513 (.A(_1217_),
    .X(net513),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout514 (.A(net516),
    .X(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout515 (.A(net516),
    .X(net515),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout516 (.A(_1231_),
    .X(net516),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout517 (.A(net518),
    .X(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout518 (.A(_1231_),
    .X(net518),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout519 (.A(net522),
    .X(net519),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout520 (.A(net522),
    .X(net520),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout521 (.A(net522),
    .X(net521),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout522 (.A(_1230_),
    .X(net522),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout523 (.A(net526),
    .X(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout524 (.A(net526),
    .X(net524),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout525 (.A(net526),
    .X(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout526 (.A(_1229_),
    .X(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout527 (.A(net982),
    .X(net527),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout528 (.A(net961),
    .X(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout529 (.A(net933),
    .X(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout530 (.A(net983),
    .X(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout531 (.A(net532),
    .X(net531),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout532 (.A(net986),
    .X(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout533 (.A(net978),
    .X(net533),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout534 (.A(\controller.inst_mem.addr[1] ),
    .X(net534),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout535 (.A(net536),
    .X(net535),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout536 (.A(net985),
    .X(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout537 (.A(net542),
    .X(net537),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout538 (.A(net542),
    .X(net538),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout539 (.A(net541),
    .X(net539),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout540 (.A(net541),
    .X(net540),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout541 (.A(net542),
    .X(net541),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout542 (.A(_0502_),
    .X(net542),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout543 (.A(net545),
    .X(net543),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout544 (.A(net545),
    .X(net544),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout545 (.A(_0502_),
    .X(net545),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout546 (.A(net547),
    .X(net546),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout547 (.A(net554),
    .X(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout548 (.A(net549),
    .X(net548),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout549 (.A(net550),
    .X(net549),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout550 (.A(net553),
    .X(net550),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout551 (.A(net553),
    .X(net551),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout554 (.A(net568),
    .X(net554),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout555 (.A(net557),
    .X(net555),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout556 (.A(net557),
    .X(net556),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout557 (.A(net558),
    .X(net557),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout558 (.A(net568),
    .X(net558),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout559 (.A(net561),
    .X(net559),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout560 (.A(net561),
    .X(net560),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout561 (.A(net568),
    .X(net561),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout562 (.A(net564),
    .X(net562),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout563 (.A(net564),
    .X(net563),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout564 (.A(net567),
    .X(net564),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout565 (.A(net567),
    .X(net565),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout566 (.A(net567),
    .X(net566),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout567 (.A(net568),
    .X(net567),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout568 (.A(net624),
    .X(net568),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout569 (.A(net570),
    .X(net569),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout570 (.A(net571),
    .X(net570),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout571 (.A(net580),
    .X(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout572 (.A(net574),
    .X(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout573 (.A(net574),
    .X(net573),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout574 (.A(net579),
    .X(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout575 (.A(net579),
    .X(net575),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout576 (.A(net578),
    .X(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout577 (.A(net579),
    .X(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout578 (.A(net579),
    .X(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout580 (.A(net624),
    .X(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout581 (.A(net584),
    .X(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout582 (.A(net584),
    .X(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout583 (.A(net584),
    .X(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout584 (.A(net591),
    .X(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout585 (.A(net586),
    .X(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout586 (.A(net587),
    .X(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout587 (.A(net591),
    .X(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout588 (.A(net589),
    .X(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout589 (.A(net591),
    .X(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout590 (.A(net591),
    .X(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout591 (.A(net605),
    .X(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout592 (.A(net594),
    .X(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout593 (.A(net594),
    .X(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout594 (.A(net605),
    .X(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout595 (.A(net596),
    .X(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout596 (.A(net597),
    .X(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout597 (.A(net605),
    .X(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout598 (.A(net604),
    .X(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout599 (.A(net603),
    .X(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout600 (.A(net603),
    .X(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout601 (.A(net602),
    .X(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout603 (.A(net604),
    .X(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout604 (.A(net605),
    .X(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout605 (.A(net624),
    .X(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout606 (.A(net607),
    .X(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout607 (.A(net623),
    .X(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout608 (.A(net611),
    .X(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout609 (.A(net610),
    .X(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout610 (.A(net611),
    .X(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout611 (.A(net623),
    .X(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout612 (.A(net614),
    .X(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout613 (.A(net614),
    .X(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout614 (.A(net623),
    .X(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout615 (.A(net616),
    .X(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout616 (.A(net622),
    .X(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout617 (.A(net622),
    .X(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout618 (.A(net622),
    .X(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout619 (.A(net621),
    .X(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout620 (.A(net621),
    .X(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout624 (.A(_1309_),
    .X(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout625 (.A(net626),
    .X(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout626 (.A(net627),
    .X(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout627 (.A(net635),
    .X(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout628 (.A(net629),
    .X(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout629 (.A(net631),
    .X(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout630 (.A(net631),
    .X(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout631 (.A(net635),
    .X(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout632 (.A(net634),
    .X(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout633 (.A(net634),
    .X(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout635 (.A(net663),
    .X(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout636 (.A(net637),
    .X(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout637 (.A(net663),
    .X(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout639 (.A(net641),
    .X(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout640 (.A(net641),
    .X(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout641 (.A(net663),
    .X(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout642 (.A(net645),
    .X(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout643 (.A(net645),
    .X(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout645 (.A(net654),
    .X(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout646 (.A(net654),
    .X(net646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout647 (.A(net654),
    .X(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout648 (.A(net650),
    .X(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout649 (.A(net650),
    .X(net649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout650 (.A(net654),
    .X(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout651 (.A(net652),
    .X(net651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout652 (.A(net653),
    .X(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout653 (.A(net654),
    .X(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout654 (.A(net663),
    .X(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout655 (.A(net657),
    .X(net655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout656 (.A(net657),
    .X(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout657 (.A(net659),
    .X(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout658 (.A(net659),
    .X(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout659 (.A(net663),
    .X(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout660 (.A(net662),
    .X(net660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout661 (.A(net662),
    .X(net661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout662 (.A(net663),
    .X(net662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout663 (.A(rst_n),
    .X(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(uio_in[7]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_can_lehmann_fsm_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net23));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_leaf_2_clk),
    .VSS(VGND));
 sg13g2_inv_8 clkload1 (.A(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_leaf_7_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_leaf_13_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload8 (.VDD(VPWR),
    .A(clknet_leaf_32_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload11 (.VDD(VPWR),
    .A(clknet_leaf_22_clk),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\controller.inst_mem.mem_data[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0273_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold3 (.A(\controller.inst_mem.mem_data[141] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold5 (.A(\controller.inst_mem.mem_data[144] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0064_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold7 (.A(\controller.inst_mem.extended_word[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0124_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold9 (.A(\controller.inst_mem.mem_data[168] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0088_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold11 (.A(\controller.inst_mem.mem_data[161] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0081_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold13 (.A(\controller.inst_mem.mem_data[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold15 (.A(\controller.inst_mem.mem_data[93] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold17 (.A(\controller.const_data[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0228_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold19 (.A(\controller.inst_mem.mem_data[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0282_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold21 (.A(\controller.const_data[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0224_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold23 (.A(\controller.inst_mem.mem_data[167] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold24 (.A(\controller.inst_mem.mem_data[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold26 (.A(\controller.inst_mem.extended_word[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold28 (.A(\controller.inst_mem.mem_data[138] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0058_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold30 (.A(\controller.inst_mem.mem_data[150] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0070_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold32 (.A(\controller.inst_mem.mem_data[165] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0085_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold34 (.A(\controller.inst_mem.mem_data[149] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold35 (.A(\controller.inst_mem.mem_data[122] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold37 (.A(\controller.inst_mem.extended_word[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0138_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold39 (.A(\controller.inst_mem.mem_data[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0283_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold41 (.A(\controller.inst_mem.mem_data[142] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold43 (.A(\controller.inst_mem.mem_data[88] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold45 (.A(\controller.const_data[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0221_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold47 (.A(\controller.inst_mem.mem_data[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0274_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold49 (.A(\controller.extended_state[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0144_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold51 (.A(\controller.inst_mem.mem_data[183] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0103_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold53 (.A(\controller.inst_mem.mem_data[190] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0110_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold55 (.A(\controller.inst_mem.mem_data[125] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0045_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold57 (.A(\controller.inst_mem.mem_data[133] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold59 (.A(\controller.inst_mem.mem_data[113] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold61 (.A(\controller.inst_mem.mem_data[104] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold63 (.A(\controller.const_data[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0218_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold65 (.A(\controller.inst_mem.extended_word[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0139_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold67 (.A(\controller.inst_mem.mem_data[191] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0111_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold69 (.A(\controller.const_data[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0236_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold71 (.A(\controller.inst_mem.mem_data[180] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0100_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold73 (.A(\controller.inst_mem.mem_data[194] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold75 (.A(\controller.inst_mem.mem_data[160] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold76 (.A(\controller.inst_mem.extended_word[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0140_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold78 (.A(\controller.inst_mem.mem_data[130] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold80 (.A(\controller.inst_mem.mem_data[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0257_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold82 (.A(\controller.const_data[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold83 (.A(\controller.const_data[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold84 (.A(\controller.inst_mem.mem_data[139] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0059_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold86 (.A(\controller.inst_mem.mem_data[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold87 (.A(\controller.inst_mem.mem_data[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold89 (.A(\controller.inst_mem.mem_data[106] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold91 (.A(\controller.const_data[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold92 (.A(\controller.const_data[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0213_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold94 (.A(\controller.inst_mem.mem_data[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold96 (.A(\controller.inst_mem.mem_data[90] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold98 (.A(\controller.inst_mem.mem_data[166] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold99 (.A(\controller.inst_mem.mem_data[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0266_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold101 (.A(\controller.inst_mem.mem_data[134] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold103 (.A(\controller.inst_mem.mem_data[185] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0105_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold105 (.A(\controller.inst_mem.mem_data[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0260_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold107 (.A(\controller.inst_mem.mem_data[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold108 (.A(\controller.inst_mem.mem_data[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold109 (.A(\controller.inst_mem.mem_data[147] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0067_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold111 (.A(\controller.inst_mem.mem_data[188] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0108_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold113 (.A(\controller.const_data[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0238_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold115 (.A(\controller.inst_mem.mem_data[91] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold117 (.A(\controller.inst_mem.mem_data[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0254_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold119 (.A(\controller.inst_mem.mem_data[126] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold121 (.A(\controller.inst_mem.mem_data[135] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold122 (.A(\controller.inst_mem.mem_data[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0280_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold124 (.A(\controller.const_data[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0209_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold126 (.A(\controller.inst_mem.mem_data[116] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0036_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold128 (.A(\controller.inst_mem.mem_data[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0277_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold130 (.A(\controller.inst_mem.mem_data[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0002_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold132 (.A(\controller.inst_mem.mem_data[145] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0065_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold134 (.A(\controller.const_data[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold135 (.A(\controller.inst_mem.mem_data[193] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold136 (.A(\controller.inst_mem.extended_word[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold137 (.A(\controller.inst_mem.mem_data[92] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold138 (.A(\controller.extended_then_action[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0134_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold140 (.A(\controller.const_data[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold142 (.A(\controller.const_data[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0239_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold144 (.A(\controller.inst_mem.mem_data[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold145 (.A(\controller.inst_mem.mem_data[132] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold146 (.A(\controller.inst_mem.mem_data[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold147 (.A(\controller.const_data[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold148 (.A(\controller.const_data[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0210_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold150 (.A(\controller.inst_mem.mem_data[177] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0097_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold152 (.A(\controller.inst_mem.mem_data[175] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0095_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold154 (.A(\controller.inst_mem.extended_word[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0126_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold156 (.A(\controller.inst_mem.mem_data[155] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0075_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold158 (.A(\controller.inst_mem.mem_data[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold159 (.A(\controller.inst_mem.mem_data[179] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold160 (.A(\controller.const_data[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold161 (.A(\controller.inst_mem.mem_data[98] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold163 (.A(\controller.inst_mem.extended_word[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold164 (.A(\controller.inst_mem.mem_data[197] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0117_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold166 (.A(\controller.const_data[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold167 (.A(\controller.inst_mem.mem_data[164] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold168 (.A(\controller.const_data[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0215_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold170 (.A(\controller.inst_mem.mem_data[189] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold171 (.A(\controller.const_data[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0230_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold173 (.A(\controller.inst_mem.mem_data[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0242_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold175 (.A(\controller.inst_mem.mem_data[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0249_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold177 (.A(\controller.inst_mem.mem_data[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold179 (.A(\controller.inst_mem.mem_data[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0263_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold181 (.A(\controller.extended_then_action[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold182 (.A(\controller.inst_mem.extended_word[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold183 (.A(\controller.inst_mem.mem_data[111] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold185 (.A(\controller.inst_mem.mem_data[163] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold186 (.A(\controller.inst_mem.mem_data[178] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold187 (.A(\controller.inst_mem.mem_data[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold188 (.A(\controller.inst_mem.mem_data[148] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold189 (.A(\controller.const_data[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold190 (.A(\controller.inst_mem.mem_data[121] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold191 (.A(\controller.inst_mem.mem_data[174] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold192 (.A(\controller.inst_mem.mem_data[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold193 (.A(\controller.inst_mem.mem_data[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0251_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold195 (.A(\controller.inst_mem.mem_data[123] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold197 (.A(\controller.inst_mem.mem_data[171] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0091_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold199 (.A(\controller.inst_mem.mem_data[124] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold200 (.A(\controller.inst_mem.mem_data[140] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold201 (.A(\controller.inst_mem.mem_data[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0244_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold203 (.A(\controller.inst_mem.mem_data[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold204 (.A(\controller.extended_state[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0145_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold206 (.A(\controller.inst_mem.mem_data[169] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0089_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold208 (.A(\controller.inst_mem.mem_data[198] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0118_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold210 (.A(\controller.inst_mem.mem_data[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold211 (.A(\controller.inst_mem.mem_data[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0271_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold213 (.A(\controller.inst_mem.mem_data[120] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold214 (.A(\controller.inst_mem.extended_word[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0128_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold216 (.A(\controller.inst_mem.mem_data[114] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0034_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold218 (.A(\controller.inst_mem.mem_data[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0267_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold220 (.A(\controller.inst_mem.mem_data[67] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold221 (.A(\controller.inst_mem.mem_data[118] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0038_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold223 (.A(\controller.inst_mem.mem_data[89] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold224 (.A(\controller.inst_mem.mem_data[152] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0072_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold226 (.A(\controller.inst_mem.mem_data[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold227 (.A(\controller.const_data[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold228 (.A(\controller.inst_mem.mem_data[107] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold230 (.A(\controller.inst_mem.mem_data[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold231 (.A(\controller.inst_mem.mem_data[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold232 (.A(\controller.inst_mem.mem_data[117] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold233 (.A(\controller.inst_mem.mem_data[170] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold234 (.A(\controller.inst_mem.mem_data[143] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold235 (.A(\controller.inst_mem.extended_word[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold236 (.A(\controller.inst_mem.extended_word[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold237 (.A(\controller.inst_mem.mem_data[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold239 (.A(\controller.inst_mem.mem_data[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0261_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold241 (.A(\controller.const_data[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold242 (.A(\controller.inst_mem.mem_data[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold243 (.A(\controller.inst_mem.mem_data[195] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0115_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold245 (.A(\controller.inst_mem.mem_data[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0284_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold247 (.A(\controller.inst_mem.mem_data[158] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0078_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold249 (.A(\controller.inst_mem.mem_data[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold250 (.A(\controller.inst_mem.mem_data[151] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold251 (.A(\controller.inst_mem.mem_data[127] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold252 (.A(\controller.inst_mem.mem_data[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold253 (.A(\controller.inst_mem.mem_data[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold254 (.A(\controller.inst_mem.mem_data[94] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold256 (.A(\controller.inst_mem.mem_data[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold257 (.A(\controller.inst_mem.mem_data[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold258 (.A(\controller.inst_mem.mem_data[105] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold259 (.A(\controller.inst_mem.mem_data[146] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold260 (.A(\controller.inst_mem.mem_data[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0269_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold262 (.A(\controller.inst_mem.mem_data[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold263 (.A(\controller.inst_mem.mem_data[173] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold264 (.A(\controller.const_data[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold265 (.A(\controller.inst_mem.mem_data[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold266 (.A(\controller.inst_mem.mem_data[192] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold267 (.A(\controller.inst_mem.mem_data[186] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0106_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold269 (.A(\controller.inst_mem.mem_data[99] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold271 (.A(\controller.const_data[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold272 (.A(\controller.inst_mem.mem_data[115] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold273 (.A(\controller.const_data[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold274 (.A(\controller.inst_mem.mem_data[95] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold275 (.A(\controller.const_data[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold276 (.A(\controller.inst_mem.mem_data[154] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold277 (.A(\controller.const_data[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold278 (.A(\controller.inst_mem.mem_data[172] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold279 (.A(\controller.inst_mem.mem_data[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0286_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold281 (.A(\controller.inst_mem.mem_data[110] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold282 (.A(\controller.inst_mem.mem_data[199] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0119_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold284 (.A(\controller.inst_mem.mem_data[131] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold285 (.A(\controller.const_data[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0211_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold287 (.A(\controller.inst_mem.mem_data[187] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold288 (.A(\controller.inst_mem.mem_data[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold289 (.A(\controller.inst_mem.mem_data[100] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold291 (.A(\controller.const_data[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold292 (.A(\controller.inst_mem.mem_data[119] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold293 (.A(\controller.const_data[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold294 (.A(\controller.inst_mem.mem_data[153] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold295 (.A(\controller.extended_jump_target[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold296 (.A(\controller.inst_mem.mem_data[196] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold297 (.A(\controller.extended_jump_target[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0120_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold299 (.A(\controller.inst_mem.mem_data[184] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold300 (.A(\controller.inst_mem.mem_data[66] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold301 (.A(\controller.inst_mem.mem_data[181] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold303 (.A(\controller.inst_mem.mem_data[176] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold304 (.A(\controller.inst_mem.mem_data[162] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold305 (.A(\controller.inst_mem.mem_data[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold306 (.A(\controller.inst_mem.mem_data[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold307 (.A(\controller.extended_jump_target[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold308 (.A(\controller.inst_mem.mem_data[109] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold309 (.A(\controller.inst_mem.mem_data[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold310 (.A(\controller.inst_mem.mem_data[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold311 (.A(\controller.extended_then_action[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold312 (.A(\controller.inst_mem.mem_data[108] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold313 (.A(\controller.inst_mem.mem_data[101] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold315 (.A(\controller.inst_mem.mem_data[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold316 (.A(\controller.inst_mem.mem_data[182] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold317 (.A(\controller.inst_mem.mem_data[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold318 (.A(\controller.inst_mem.mem_data[102] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold320 (.A(\controller.inst_mem.mem_data[157] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold321 (.A(\controller.inst_mem.mem_data[103] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold322 (.A(\controller.inst_mem.mem_data[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0246_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold324 (.A(\controller.inst_mem.mem_data[159] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold325 (.A(\controller.inst_mem.mem_data[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold326 (.A(\controller.const_data[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold327 (.A(\controller.inst_mem.mem_data[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold328 (.A(\controller.inst_mem.mem_data[156] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold329 (.A(\controller.inst_mem.mem_data[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold330 (.A(\controller.inst_mem.mem_data[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold331 (.A(\controller.extended_then_action[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold332 (.A(\controller.counter2.counter_0[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold334 (.A(\controller.extended_then_action[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold335 (.A(\controller.extended_then_action[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold336 (.A(\controller.counter2.counter_1[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0203_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold338 (.A(\controller.extended_cond.opcode[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold339 (.A(\controller.counter2.counter_0[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0185_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold341 (.A(\controller.counter2.counter_1[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0198_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold343 (.A(\controller.counter2.counter_1[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0195_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold345 (.A(\controller.counter2.counter_1[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold346 (.A(\controller.counter2.counter_0[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold347 (.A(\controller.counter2.counter_0[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0182_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold349 (.A(\controller.counter2.counter_0[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold350 (.A(\controller.counter2.counter_0[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0187_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold352 (.A(\controller.counter2.counter_0[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0189_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold354 (.A(\controller.counter2.counter_1[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0201_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold356 (.A(\controller.counter2.counter_1[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold357 (.A(\controller.counter2.counter_1[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold359 (.A(\controller.counter2.counter_0[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold360 (.A(\controller.counter2.counter_1[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0202_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold362 (.A(\controller.counter2.counter_1[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold363 (.A(\controller.counter2.counter_1[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold364 (.A(\controller.counter2.counter_1[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0194_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold366 (.A(\controller.alu_buffer.buffer[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0172_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold368 (.A(\controller.counter2.counter_1[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold369 (.A(\controller.counter2.counter_0[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold370 (.A(\controller.output_controller.keep[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0175_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold372 (.A(\controller.counter2.counter_0[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0178_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold374 (.A(\controller.counter2.counter_1[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold375 (.A(\controller.alu_buffer.buffer[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold377 (.A(\controller.counter2.counter_0[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0186_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold379 (.A(\controller.counter2.counter_1[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0205_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold381 (.A(\controller.counter2.counter_0[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0179_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold383 (.A(\controller.counter2.counter_0[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold385 (.A(\controller.counter2.counter_1[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold386 (.A(\controller.alu_buffer.buffer[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0644_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0159_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold389 (.A(\controller.extended_cond.opcode[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0129_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold391 (.A(\controller.counter2.counter_0[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold393 (.A(\controller.output_controller.keep[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0174_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold395 (.A(\controller.counter2.counter_1[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold396 (.A(\controller.extended_cond.opcode[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold397 (.A(\controller.counter2.counter_0[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold398 (.A(\controller.alu_buffer.buffer[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0168_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold400 (.A(\controller.counter2.counter_0[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold401 (.A(\controller.alu_buffer.buffer[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0169_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold403 (.A(\controller.alu_buffer.buffer[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0163_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold405 (.A(\controller.alu_buffer.buffer[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0167_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold407 (.A(\controller.alu_buffer.buffer[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0162_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold409 (.A(\controller.alu_buffer.buffer[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0171_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold411 (.A(\controller.alu_buffer.buffer[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0166_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold413 (.A(\controller.alu_buffer.buffer[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold414 (.A(\controller.alu_buffer.buffer[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0155_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold416 (.A(\controller.alu_buffer.buffer[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0158_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold418 (.A(\controller.alu_buffer.buffer[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0165_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold420 (.A(\controller.alu_buffer.buffer[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0149_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold422 (.A(\controller.alu_buffer.buffer[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0161_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold424 (.A(\controller.alu_buffer.buffer[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0150_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold426 (.A(\controller.alu_buffer.buffer[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold428 (.A(\controller.alu_buffer.buffer[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0160_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold430 (.A(\controller.alu_buffer.buffer[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold431 (.A(\controller.inst_mem.addr[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0147_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold433 (.A(\controller.alu_buffer.buffer[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0154_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold435 (.A(\controller.alu_buffer.buffer[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold436 (.A(\controller.alu_buffer.buffer[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold437 (.A(\controller.alu_buffer.buffer[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold438 (.A(\controller.inst_mem.addr[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold439 (.A(\controller.inst_mem.addr[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0148_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net987));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(ui_in[0]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(ui_in[2]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(ui_in[3]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(ui_in[5]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(ui_in[6]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[0]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[1]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[2]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[4]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[5]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[6]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[7]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(ui_in[1]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(uio_in[3]));
 sg13g2_fill_2 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_501 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net23;
 assign uio_oe[1] = net24;
 assign uio_oe[2] = net25;
 assign uio_oe[3] = net26;
 assign uio_oe[4] = net27;
 assign uio_oe[5] = net28;
 assign uio_oe[6] = net29;
 assign uio_oe[7] = net30;
 assign uio_out[0] = net31;
 assign uio_out[1] = net32;
 assign uio_out[2] = net33;
 assign uio_out[3] = net34;
 assign uio_out[4] = net35;
 assign uio_out[5] = net36;
 assign uio_out[6] = net37;
 assign uio_out[7] = net38;
endmodule
